library ieee;
use ieee.std_logic_1164.all;
use work.Common.all;

entity test_conv2d is
	port (
	 clk : in std_logic;
	 filtered_img : out img_1d_vec_float (0 to (row*col) - 1) := (others => (others => '0'))
	);
end entity;

architecture rch of test_conv2d is
	
	component conv2d is
	generic (
		row : integer := 10;
		col : integer := 10;
		m : integer := 7;
		n : integer := 7
	);
	port (
		clk : in std_logic;
		img : in img_1d_vec_float (0 to (row*col) - 1);
		mask : in img_1d_vec_float(0 to (m*n) - 1);
		filtered_img : out img_1d_vec_float (0 to (row*col) - 1) := (others => (others => '0'));
		conv2d_ready : out std_logic
	);
	end component;
	
	constant img_rom : img_1d_vec_float (0 to (row*col) - 1) := (
		"0101100111100000", "0101100111101000", "0101100111110000", "0101100111111000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101000111000", "0101101000111000", "0101101001001000", "0101101000111000", "0101101001000000", "0101101000111000", "0101101000101000", "0101101001010000", "0101101000100000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000111000", "0101101001000000", "0101101000101000", "0101101001010000", "0101101001000000", "0101101000101000", "0101101001100000", "0101101000100000", "0101101001010000", "0101101001000000", "0101101000101000", "0101101000110000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000011000", "0101101000110000", "0101101000101000", "0101101000001000", "0101101001010000", "0101101000010000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111100000", "0101100111101000", "0101100111100000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100110111000", "0101100110111000", "0101100110101000", "0101100110100000", "0101100110010000", "0101100110001000", "0101100101111000", "0101100101110000", "0101100101101000", "0101101101100000", "0101100111101000", "0101100111110000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101001001000", "0101101001001000", "0101101001000000", "0101101000011000", "0101101001011000", "0101101001010000", "0101101000100000", "0101101001010000", "0101101001000000", "0101101000100000", "0101101001100000", "0101101001001000", "0101101000110000", "0101101001010000", "0101101000101000", "0101101001001000", "0101101001100000", "0101101000111000", "0101101001001000", "0101101000100000", "0101101000111000", "0101101001011000", "0101101000101000", "0101101000111000", "0101101000011000", "0101101000111000", "0101101001000000", "0101101000110000", "0101101000101000", "0101101000110000", "0101100111111000", "0101101001000000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110111000", "0101100110110000", "0101100110101000", "0101100110011000", "0101100110010000", "0101100110001000", "0101100110001000", "0101100101111000", "0101101101101000", "0101100111110000", "0101100111110000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000000000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101001010000", "0101101000111000", "0101101001111000", "0101101001001000", "0101101000110000", "0101101001001000", "0101101000110000", "0101101000110000", "0101101001011000", "0101101000101000", "0101101000011000", "0101101001000000", "0101100110010000", "0101100111101000", "0101101001110000", "0101101001000000", "0101101000101000", "0101101001010000", "0101101001100000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000111000", "0101101000100000", "0101101001001000", "0101101000011000", "0101101000100000", "0101101000110000", "0101101000110000", "0101101001001000", "0101101000010000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111010000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110111000", "0101100110111000", "0101100110110000", "0101100110101000", "0101100110100000", "0101100110010000", "0101100110001000", "0101100101111000", "0101101101100000", "0101100111101000", "0101100111110000", "0101100111111000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000000000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101000101000", "0101101000101000", "0101001000100000", "0101010011110000", "0101100111000000", "0101000100100000", "0101011111100000", "0101100001100000", "0101100111110000", "0100101110000000", "0101100010101000", "0101010011100000", "0101100011001000", "0101101000111000", "0101101001001000", "0101101001001000", "0101101000101000", "0101101000111000", "0101101000101000", "0101101001000000", "0101101000110000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110111000", "0101100110110000", "0101100110101000", "0101100110001000", "0101100110001000", "0101100101110000", "0101101101011000", "0101100111101000", "0101100111110000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001000000", "0101101001010000", "0101101001010000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101001001000", "0101101001011000", "0101101001000000", "0101000110100000", "0101001111100000", "0101001100100000", "0101011011100000", "0101010011110000", "0101010010110000", "0101001101000000", "0100110111000000", "0100110001000000", "0100101010000000", "0100100000000000", "0100100100000000", "0100110011000000", "0101100011110000", "0101100010010000", "0101101001010000", "0101100001000000", "0101101000001000", "0101101000010000", "0101101001101000", "0101101000110000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110110000", "0101100110101000", "0101100110011000", "0101100110010000", "0101100110000000", "0101101101100000", "0101100111110000", "0101100111111000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000110000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001000000", "0101101001010000", "0101101001101000", "0101101001001000", "0101101001001000", "0101101000110000", "0101101000011000", "0101100010111000", "0101101000111000", "0101101000110000", "0101000011000000", "0101011010100000", "0100111110000000", "0101000000000000", "0100110111000000", "0100111101000000", "0101001100000000", "0100111101000000", "0100101110000000", "0100101100000000", "0100101110000000", "0100110010000000", "0100111011000000", "0100100000000000", "0101011100100000", "0101100111001000", "0101101000110000", "0101100010101000", "0101101001101000", "0101101000100000", "0101101000111000", "0101101001001000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110110000", "0101100110110000", "0101100110101000", "0101100110101000", "0101100110001000", "0101101101101000", "0101100111111000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001001000", "0101101000101000", "0101101001001000", "0101100111111000", "0100110000000000", "0101000101100000", "0101010001110000", "0101100000101000", "0100111111000000", "0100111100000000", "0101000000000000", "0100101100000000", "0101000000000000", "0101000000100000", "0101000011100000", "0101010010010000", "0101001010100000", "0101000101000000", "0100111100000000", "0100110011000000", "0101000111100000", "0100110011000000", "0100111001000000", "0101011000010000", "0101011110100000", "0101100010001000", "0101011101100000", "0101101001010000", "0101101001001000", "0101101001011000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111100000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110110000", "0101100110110000", "0101100110110000", "0101100110010000", "0101101101100000", "0101100111111000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001010000", "0101101000011000", "0101100101101000", "0100110110000000", "0101001001100000", "0101010001110000", "0101010100000000", "0101000110000000", "0101000100000000", "0101000010100000", "0100111110000000", "0100110101000000", "0101001011100000", "0101001010100000", "0101010000010000", "0101001010100000", "0101010000110000", "0101001101100000", "0101001000000000", "0101010010100000", "0101001000000000", "0101001000100000", "0101001010000000", "0101010111010000", "0101101000010000", "0101010010010000", "0101101000000000", "0101101001001000", "0101101001000000", "0101101001001000", "0101101001001000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111101000", "0101100111101000", "0101100111101000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100110111000", "0101100110111000", "0101100110111000", "0101100110110000", "0101100110010000", "0101101101101000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000111000", "0101101001000000", "0101101001001000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101001100000", "0101101001011000", "0101101000100000", "0101100010010000", "0100110100000000", "0101010101110000", "0101000110000000", "0101001000000000", "0101001000000000", "0100110011000000", "0101000001100000", "0100110000000000", "0100111001000000", "0101010000100000", "0101010000000000", "0101010010000000", "0101010001000000", "0101010100010000", "0101010001010000", "0101000101000000", "0101010100010000", "0101001010100000", "0101001011000000", "0101010010110000", "0101010100010000", "0101011100000000", "0101011111000000", "0101100100000000", "0101100101001000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101001011000", "0101101000110000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000110000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111101000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111001000", "0101100111001000", "0101100111001000", "0101100110111000", "0101100110111000", "0101100110101000", "0101101101011000", "0101101000000000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001101000", "0101101001011000", "0101101001100000", "0101101000111000", "0101010000000000", "0101000000000000", "0101011010010000", "0100110100000000", "0100110100000000", "0101000010100000", "0101000000000000", "0100111111000000", "0100111001000000", "0100100000000000", "0100111100000000", "0101000010000000", "0101000110000000", "0101000111000000", "0101000110100000", "0101010110010000", "0101000111100000", "0100101000000000", "0101000011100000", "0101000000000000", "0100111110000000", "0101010001100000", "0101001100100000", "0101010101100000", "0101010010010000", "0101100111011000", "0101100111110000", "0101101001010000", "0101101001000000", "0101101001011000", "0101101000010000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000001000", "0101101001000000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111100000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111001000", "0101100111001000", "0101100111001000", "0101100110111000", "0101100110111000", "0101100110110000", "0101101101011000", "0101101000000000", "0101101000001000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101001000000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101000101000", "0101100111010000", "0100100110000000", "0101000011000000", "0101000010100000", "0101001010000000", "0100111011000000", "0101000100100000", "0101000100000000", "0101000001100000", "0100110111000000", "0100110001000000", "0100110100000000", "0100111111000000", "0100110100000000", "0101000010100000", "0100110011000000", "0101000101100000", "0100111110000000", "0000000000000000", "0100111001000000", "0100110111000000", "0101001101000000", "0100011100000000", "0101000010000000", "0101001011000000", "0101000111000000", "0101100101011000", "0101101000001000", "0101101001010000", "0101101001100000", "0101101001001000", "0101101001100000", "0101100111111000", "0101101000111000", "0101101001000000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111110000", "0101100111110000", "0101100111111000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110110000", "0101101101100000", "0101101000001000", "0101101000010000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000111000", "0101101001001000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001001000", "0101101001011000", "0101101001000000", "0101010010010000", "0100110101000000", "0101000000000000", "0100111101000000", "0101000110000000", "0101001101100000", "0101000100000000", "0101000100000000", "0101000010000000", "0100111011000000", "0101000000000000", "0100011000000000", "0100110001000000", "0100101100000000", "0100111101000000", "0100101100000000", "0101000001000000", "0100101100000000", "0100111100000000", "0100110000000000", "0100101110000000", "0100101110000000", "0100101100000000", "0100110111000000", "0101000010100000", "0101000101000000", "0101011101110000", "0101100011101000", "0101100111010000", "0101100110111000", "0101101000110000", "0101101000010000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101001001000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111101000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110111000", "0101101101100000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101001000000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001100000", "0101101001010000", "0101000000000000", "0100111110000000", "0100111100000000", "0100111000000000", "0101000110000000", "0101001101100000", "0100110111000000", "0100101000000000", "0101000110000000", "0100101110000000", "0100110001000000", "0100101010000000", "0101001001000000", "0100110110000000", "0100110011000000", "0100110001000000", "0101001010000000", "0100111000000000", "0100110001000000", "0100111111000000", "0100110001000000", "0100110101000000", "0100110101000000", "0100101010000000", "0100110010000000", "0100110000000000", "0100110101000000", "0101011010010000", "0101011100100000", "0101010101110000", "0101001011000000", "0101001101000000", "0101010110010000", "0101101000000000", "0101101000101000", "0101101001001000", "0101101000100000", "0101101001000000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100111001000", "0101100110111000", "0101101101100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101001010000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001000000", "0101101001111000", "0100110111000000", "0101010011010000", "0100110010000000", "0100100100000000", "0100110010000000", "0100111000000000", "0100111111000000", "0101000011000000", "0100101110000000", "0101000001100000", "0100110111000000", "0100110110000000", "0100111100000000", "0100111110000000", "0100111001000000", "0101000110000000", "0101000000000000", "0101000110100000", "0101000000000000", "0101000001000000", "0101000001000000", "0100110101000000", "0100110110000000", "0100100100000000", "0100110000000000", "0100111010000000", "0101000000000000", "0100111110000000", "0101000011100000", "0101010101000000", "0101011001010000", "0101010110000000", "0101011100010000", "0101100111011000", "0101100111100000", "0101101001000000", "0101101001011000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000001000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101000001000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101100110111000", "0101101101100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000101000", "0101101000111000", "0101101001001000", "0101101001011000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101011110100000", "0100110000000000", "0100111010000000", "0100110100000000", "0100110010000000", "0100100110000000", "0100110010000000", "0100101100000000", "0100111101000000", "0101000100000000", "0101000111000000", "0101000100000000", "0101001001000000", "0101000110000000", "0101001001000000", "0101010110000000", "0101011000010000", "0101010110110000", "0101010101110000", "0101010101010000", "0101010100010000", "0101001010100000", "0101000100100000", "0100101110000000", "0100101100000000", "0100011100000000", "0101000111100000", "0100101000000000", "0101000100100000", "0101001111000000", "0101001110100000", "0101010010100000", "0101100010011000", "0101100001000000", "0101101000010000", "0101101001101000", "0101101000111000", "0101101001000000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000001000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111010000", "0101100111001000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100110111000", "0101101101101000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000101000", "0101101000111000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001000000", "0101100100111000", "0100110110000000", "0100101110000000", "0100101100000000", "0100100100000000", "0100100110000000", "0100101000000000", "0100110000000000", "0101000100100000", "0101010100110000", "0101010011000000", "0101010101000000", "0101010111010000", "0101011100000000", "0101011111010000", "0101100011101000", "0101100110001000", "0101100011100000", "0101100111001000", "0101101001101000", "0101100110111000", "0101100010110000", "0101100110000000", "0101010111010000", "0101010000110000", "0100110111000000", "0100101010000000", "0100100100000000", "0100101100000000", "0101000000000000", "0100110111000000", "0101000010100000", "0101010001010000", "0101010011110000", "0101100100111000", "0101101001001000", "0101101000100000", "0101101001100000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111001000", "0101100111001000", "0101100111000000", "0101100111000000", "0101100111000000", "0101101101101000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000101000", "0101101000110000", "0101101001010000", "0101101001100000", "0101101001011000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001111000", "0101101001100000", "0101101001000000", "0101101001101000", "0101101000011000", "0101100111011000", "0101101000100000", "0101100111110000", "0100110101000000", "0100101100000000", "0100101010000000", "0100101010000000", "0100010000000000", "0100101110000000", "0100100000000000", "0101000101000000", "0101010101110000", "0101011111100000", "0101100000000000", "0101100011101000", "0101100110000000", "0101100111010000", "0101101000100000", "0101101011000000", "0101101100000000", "0101101011111000", "0101101101001000", "0101101101000000", "0101101100101000", "0101101100101000", "0101101100000000", "0101101001001000", "0101100010110000", "0101000000000000", "0100101010000000", "0100011000000000", "0101001110000000", "0101001101100000", "0101010010000000", "0101001000100000", "0101001110100000", "0101010011110000", "0101100011110000", "0101100101001000", "0101101000000000", "0101101001000000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111010000", "0101100111000000", "0101100111000000", "0101100111001000", "0101100111000000", "0101101101100000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000111000", "0101101001000000", "0101101001011000", "0101101001011000", "0101101001001000", "0101101001100000", "0101101001100000", "0101101010000000", "0101101001000000", "0101101001100000", "0101101001101000", "0101101001010000", "0101101001001000", "0101100100111000", "0101011010110000", "0101011001010000", "0100100100000000", "0100011100000000", "0100100000000000", "0100011000000000", "0011110000000000", "0100101110000000", "0101000101100000", "0101010110010000", "0101100000000000", "0101100100001000", "0101100110101000", "0101100111111000", "0101101001111000", "0101101010001000", "0101101011110000", "0101101100101000", "0101101101001000", "0101101100110000", "0101101101010000", "0101101101000000", "0101101100100000", "0101101100011000", "0101101011111000", "0101101011011000", "0101101010011000", "0101011001100000", "0100111111000000", "0100110000000000", "0101000001000000", "0100100010000000", "0101000110000000", "0101001001100000", "0101010000000000", "0101011001010000", "0101011000010000", "0101101000111000", "0101101001011000", "0101101001001000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111001000", "0101100111000000", "0101101101100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101001001000", "0101101001010000", "0101101001100000", "0101101001011000", "0101101001000000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001010000", "0101101001011000", "0101101001101000", "0101101010001000", "0101101000111000", "0101101000110000", "0101100000101000", "0101011010010000", "0100110000000000", "0100100110000000", "0100000000000000", "0100011100000000", "0100000000000000", "0101001000000000", "0101010100010000", "0101011110000000", "0101100010101000", "0101100110001000", "0101101000000000", "0101101001100000", "0101101010101000", "0101101100001000", "0101101100101000", "0101101100100000", "0101101100100000", "0101101100101000", "0101101100011000", "0101101100100000", "0101101100010000", "0101101100010000", "0101101100000000", "0101101011101000", "0101101011011000", "0101100101000000", "0101000010000000", "0100100110000000", "0101000101100000", "0101001110100000", "0101001010100000", "0101000101000000", "0101001000100000", "0100101110000000", "0101100101010000", "0101100111011000", "0101101000110000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111010000", "0101100111001000", "0101100111000000", "0101100111001000", "0101100110111000", "0101101101100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101001001000", "0101101001010000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001100000", "0101101001101000", "0101101001010000", "0101101001111000", "0101101001101000", "0101101001011000", "0101101000110000", "0101101001100000", "0101101001011000", "0101101000100000", "0101011111000000", "0100111100000000", "0100110000000000", "0100010100000000", "0000000000000000", "0100011100000000", "0101010011000000", "0101011101000000", "0101100010001000", "0101100101011000", "0101100111100000", "0101101001011000", "0101101010110000", "0101101011100000", "0101101100100000", "0101101100011000", "0101101100110000", "0101101100100000", "0101101100111000", "0101101100010000", "0101101100100000", "0101101100001000", "0101101100000000", "0101101011111000", "0101101011110000", "0101101010101000", "0101101011010000", "0101010011110000", "0100111010000000", "0100110110000000", "0101000101100000", "0101010000110000", "0101000000100000", "0100110001000000", "0101000001100000", "0101000110000000", "0101101000110000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111001000", "0101100111001000", "0101100111000000", "0101101101100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000101000", "0101101000111000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001001000", "0101101001101000", "0101101001110000", "0101101001011000", "0101101001101000", "0101101001011000", "0101101001110000", "0101101001100000", "0101101001110000", "0101101001001000", "0101101000100000", "0101000110000000", "0101001011000000", "0100100110000000", "0100011100000000", "0100010000000000", "0100111101000000", "0101010101000000", "0101100000100000", "0101100011111000", "0101100110010000", "0101101000100000", "0101101001000000", "0101101011111000", "0101101010100000", "0101101100010000", "0101101100010000", "0101101100101000", "0101101100101000", "0101101101010000", "0101101100101000", "0101101100111000", "0101101100011000", "0101101100000000", "0101101011101000", "0101101011011000", "0101101100000000", "0101101010111000", "0101100010100000", "0101000011000000", "0100101010000000", "0100110110000000", "0100111110000000", "0101001000000000", "0101001001100000", "0101000000000000", "0101010101110000", "0101101000000000", "0101101001000000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111100000", "0101100111011000", "0101100111001000", "0101100111010000", "0101100111000000", "0101101101100000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000010000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000111000", "0101101001001000", "0101101001010000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001000000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001011000", "0101101001111000", "0101011111010000", "0101001001000000", "0100111110000000", "0100001000000000", "0000000000000000", "0100100010000000", "0101001101000000", "0101011010010000", "0101100001011000", "0101100100000000", "0101100111101000", "0101101000011000", "0101101001110000", "0101101010010000", "0101101011001000", "0101101011110000", "0101101100101000", "0101101011110000", "0101101100010000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101100101000", "0101101100011000", "0101101011110000", "0101101011100000", "0101101010001000", "0101101001100000", "0101100011011000", "0101010110110000", "0100100110000000", "0101000100000000", "0100110001000000", "0101000000000000", "0100111101000000", "0101001010000000", "0101011011010000", "0101101001011000", "0101101001001000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111100000", "0101100111011000", "0101100111010000", "0101100111010000", "0101100111000000", "0101101101100000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000110000", "0101101000101000", "0101101001000000", "0101101001010000", "0101101001001000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001111000", "0101101001111000", "0101101001101000", "0101101001100000", "0101100111001000", "0100101010000000", "0100110001000000", "0100010100000000", "0100110001000000", "0101010011110000", "0101011101110000", "0101100001111000", "0101100100010000", "0101100111110000", "0101101001011000", "0101101010010000", "0101101010011000", "0101101011100000", "0101101100000000", "0101101011110000", "0101101011111000", "0101101100101000", "0101101100100000", "0101101100111000", "0101101100101000", "0101101100100000", "0101101100100000", "0101101011111000", "0101101011010000", "0101101011001000", "0101101010011000", "0101100111000000", "0101010110100000", "0101000100100000", "0100101000000000", "0100101110000000", "0101000000100000", "0101000101100000", "0101010000000000", "0101100101001000", "0101101001010000", "0101101001100000", "0101101001010000", "0101101001110000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111011000", "0101100111011000", "0101100111001000", "0101101101101000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101001010000", "0101101001011000", "0101101001001000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001111000", "0101100111100000", "0101000100000000", "0100010000000000", "0100011000000000", "0101000101100000", "0101010111010000", "0101011110100000", "0101100010010000", "0101100100111000", "0101100110111000", "0101101000001000", "0101101010001000", "0101101001111000", "0101101011101000", "0101101100010000", "0101101100011000", "0101101011100000", "0101101100100000", "0101101011111000", "0101101100100000", "0101101100010000", "0101101100011000", "0101101100101000", "0101101100000000", "0101101011010000", "0101101011000000", "0101101010100000", "0101100111110000", "0101011101010000", "0101001100000000", "0100100110000000", "0100010000000000", "0100101010000000", "0100101010000000", "0100110011000000", "0101101000001000", "0101101000101000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101000110000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111100000", "0101100111001000", "0101101101101000", "0101101000011000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001101000", "0100100010000000", "0100001000000000", "0100110000000000", "0101001010100000", "0101011001100000", "0101100000001000", "0101100010110000", "0101100101111000", "0101100101101000", "0101101000100000", "0101101001010000", "0101101010101000", "0101101100000000", "0101101100000000", "0101101011101000", "0101101011111000", "0101101100011000", "0101101100010000", "0101101100010000", "0101101100000000", "0101101100110000", "0101101100101000", "0101101100110000", "0101101100001000", "0101101011111000", "0101101010110000", "0101100100111000", "0101011110110000", "0101010010010000", "0100111010000000", "0100101010000000", "0100110100000000", "0100110110000000", "0100110111000000", "0101101001111000", "0101101001100000", "0101101001010000", "0101101001101000", "0101101001101000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111100000", "0101101101011000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101001001000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101010001000", "0100110010000000", "0100101100000000", "0100110010000000", "0101001100000000", "0101011100010000", "0101011111110000", "0101100010010000", "0101100011110000", "0101100101011000", "0101100111101000", "0101101000110000", "0101101010101000", "0101101100010000", "0101101100110000", "0101101100001000", "0101101011101000", "0101101101001000", "0101101100000000", "0101101100010000", "0101101100011000", "0101101100010000", "0101101100100000", "0101101101100000", "0101101100111000", "0101101011110000", "0101101010111000", "0101100110010000", "0101100000010000", "0101001101000000", "0100110101000000", "0100101100000000", "0100110011000000", "0101000001000000", "0101000110100000", "0101101000111000", "0101101001110000", "0101101001110000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101100111100000", "0101101101011000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101000111000", "0101101001000000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000111000", "0101101001000000", "0101101001000000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101010000000", "0101010100100000", "0100110010000000", "0100111000000000", "0101010011100000", "0101011100100000", "0101100001001000", "0101100100001000", "0101100100100000", "0101100110101000", "0101100111110000", "0101101001110000", "0101101011100000", "0101101100011000", "0101101100100000", "0101101100011000", "0101101100010000", "0101101100100000", "0101101101010000", "0101101100101000", "0101101100111000", "0101101100011000", "0101101100101000", "0101101100101000", "0101101101010000", "0101101100001000", "0101101011010000", "0101100110100000", "0101011100110000", "0101010010100000", "0100101010000000", "0100100100000000", "0100111101000000", "0100110010000000", "0101001010000000", "0101101000001000", "0101101001110000", "0101101010000000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111101000", "0101100111100000", "0101101101011000", "0101101000101000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001001000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010011000", "0101100100100000", "0100100110000000", "0100111001000000", "0101011001110000", "0101011101010000", "0101100001101000", "0101100010110000", "0101100011111000", "0101100110100000", "0101101000010000", "0101101011000000", "0101101100001000", "0101101100101000", "0101101011111000", "0101101011110000", "0101101011101000", "0101101101001000", "0101101101010000", "0101101101011000", "0101101101000000", "0101101101000000", "0101101100111000", "0101101101000000", "0101101011111000", "0101101100110000", "0101101010110000", "0101101000110000", "0101011010000000", "0101000001000000", "0100111111000000", "0100111000000000", "0100110010000000", "0100110011000000", "0101011100010000", "0101101010001000", "0101101001000000", "0101101001010000", "0101101010001000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111101000", "0101100111101000", "0101101101100000", "0101101000100000", "0101101000110000", "0101101000111000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010010000", "0101101001100000", "0100110100000000", "0101000001000000", "0101011001000000", "0101011110000000", "0101100010001000", "0101100011101000", "0101100100110000", "0101100111011000", "0101101001111000", "0101101011100000", "0101101011100000", "0101101101001000", "0101101100011000", "0101101100011000", "0101101100100000", "0101101100110000", "0101101101010000", "0101101101101000", "0101101101010000", "0101101101100000", "0101101101011000", "0101101100011000", "0101101100101000", "0101101100010000", "0101101010110000", "0101101100000000", "0101100111100000", "0101011001000000", "0101001001000000", "0101000010100000", "0100100110000000", "0100100100000000", "0101100011110000", "0101101001111000", "0101101010000000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111110000", "0101100111110000", "0101101101100000", "0101101000101000", "0101101000110000", "0101101001000000", "0101101001000000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010000000", "0100110011000000", "0101001010000000", "0101011010000000", "0101011110000000", "0101100001101000", "0101100011011000", "0101100101100000", "0101100111000000", "0101101001110000", "0101101011000000", "0101101010111000", "0101101100110000", "0101101011110000", "0101101100010000", "0101101100010000", "0101101101000000", "0101101110000000", "0101101110011000", "0101101101111000", "0101101110000000", "0101101100111000", "0101101101101000", "0101101011110000", "0101101100100000", "0101101010110000", "0101101010100000", "0101101010011000", "0101100000010000", "0101001010100000", "0101000101100000", "0100101010000000", "0100111010000000", "0101101001010000", "0101101001001000", "0101101001100000", "0101101010001000", "0101101001111000", "0101101001011000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111110000", "0101100111110000", "0101101101100000", "0101101000110000", "0101101001000000", "0101101001001000", "0101101001010000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010100000", "0100101100000000", "0101001110100000", "0101011001100000", "0101011100100000", "0101100011010000", "0101100011111000", "0101100110110000", "0101101000000000", "0101101010000000", "0101101010010000", "0101101010010000", "0101101011101000", "0101101011010000", "0101101101011000", "0101101101011000", "0101101100011000", "0101101101101000", "0101101101000000", "0101101100000000", "0101101010010000", "0101100100110000", "0101101100110000", "0101101100011000", "0101101010101000", "0101101011001000", "0101101010001000", "0101101010111000", "0101100100000000", "0101010110000000", "0101000110000000", "0100101110000000", "0101001011000000", "0101101001101000", "0101101010001000", "0101101010000000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111110000", "0101100111101000", "0101101101011000", "0101101000111000", "0101101001001000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001111000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010011000", "0101101010011000", "0100101010000000", "0101010000010000", "0101011001000000", "0101011011110000", "0101100000111000", "0101010101010000", "0101011010110000", "0101100010100000", "0101100111100000", "0101101001000000", "0101101001110000", "0101101010101000", "0101101001111000", "0101101011111000", "0101101010111000", "0101101011101000", "0101100100001000", "0101011000100000", "0101011011010000", "0101011110110000", "0101100111011000", "0101100011010000", "0101101010010000", "0101101011000000", "0101101011010000", "0101101010011000", "0101101001111000", "0101100110111000", "0101010011100000", "0100101110000000", "0100111110000000", "0101011101010000", "0101101010000000", "0101101010010000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101101000000000", "0101100111110000", "0101100111101000", "0101101101011000", "0101101000110000", "0101101001010000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001101000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010110000", "0101101010100000", "0100111000000000", "0101001100100000", "0101011000000000", "0101010110110000", "0101010101110000", "0101010110110000", "0101001111000000", "0101010001100000", "0101011010110000", "0101100011111000", "0101100111111000", "0101101010100000", "0101101001111000", "0101101011110000", "0101101001100000", "0101101001000000", "0101011111100000", "0101011001110000", "0101011101010000", "0101100100110000", "0101100011101000", "0101100010000000", "0101101000000000", "0101101001000000", "0101101010110000", "0101101010110000", "0101101000101000", "0101100111111000", "0101010001010000", "0101010000100000", "0101000010100000", "0101100000011000", "0101101001110000", "0101101010010000", "0101101001110000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000001000", "0101100111111000", "0101101000000000", "0101100111111000", "0101100111110000", "0101101101100000", "0101101001000000", "0101101001011000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001110000", "0101101001111000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0100111010000000", "0101001000000000", "0101011000110000", "0101010100000000", "0101011001100000", "0101011101100000", "0101100001011000", "0101011111100000", "0101011101110000", "0101011011010000", "0101100011110000", "0101100111000000", "0101101001110000", "0101101011111000", "0101101000011000", "0101100111000000", "0101100110001000", "0101100110110000", "0101101011101000", "0101101101010000", "0101101010000000", "0101101001100000", "0101100111100000", "0101101010100000", "0101101010111000", "0101101010101000", "0101101001000000", "0101100111000000", "0101010000100000", "0101010110100000", "0101010010000000", "0101011000000000", "0101101010011000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101001100000", "0101101010001000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111110000", "0101100111110000", "0101101101011000", "0101101001010000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101010000000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101011000000", "0101101010110000", "0101000101100000", "0101001000000000", "0101011000100000", "0101010110010000", "0101011000010000", "0101100001100000", "0101100101001000", "0101101001000000", "0101101011000000", "0101100110011000", "0101010110010000", "0101100011111000", "0101101010000000", "0101101101011000", "0101101010001000", "0101100101111000", "0101100111001000", "0101100010000000", "0101100001011000", "0101100100000000", "0101101100000000", "0101101010101000", "0101101000001000", "0101101001100000", "0101101010111000", "0101101010010000", "0101101000010000", "0101100110111000", "0101001011000000", "0101010110000000", "0101010110010000", "0101001110000000", "0101101010000000", "0101101010100000", "0101101001110000", "0101101010000000", "0101101010011000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111110000", "0101100111110000", "0101101101100000", "0101101001011000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101010110000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010100000", "0101010011010000", "0101000001000000", "0101011001100000", "0101011000110000", "0101010101000000", "0101100010000000", "0101100000111000", "0101100010010000", "0101101000011000", "0101011000000000", "0101011011010000", "0101011111010000", "0101101011101000", "0101101110100000", "0101101100110000", "0101100010111000", "0101011011000000", "0101010011110000", "0100111010000000", "0101011000000000", "0101100000100000", "0101101000100000", "0101101000011000", "0101101001111000", "0101101010110000", "0101101010001000", "0101101000001000", "0101100110100000", "0101010001000000", "0101011011000000", "0101011000110000", "0101011110100000", "0101101010101000", "0101101010000000", "0101101010010000", "0101101001110000", "0101101010011000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001001000", "0101101001001000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101101101000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010101000", "0101101011100000", "0101100010001000", "0100111100000000", "0101010110100000", "0101011000100000", "0101010111110000", "0101010011110000", "0101011111000000", "0101000101000000", "0101010100100000", "0101010110110000", "0101011000100000", "0101011000000000", "0101101011000000", "0101101110010000", "0101101100101000", "0101100011010000", "0101011101010000", "0101100111100000", "0101010111000000", "0101011101100000", "0101100110101000", "0101100001111000", "0101101010101000", "0101101011000000", "0101101001101000", "0101101010100000", "0101100111011000", "0101100100011000", "0101010010110000", "0101010101110000", "0101100101110000", "0101100100011000", "0101101010011000", "0101101010101000", "0101101010001000", "0101101011000000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101101101000", "0101101001100000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001011000", "0101101001101000", "0101101001110000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010100000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101011010000", "0101101011000000", "0101100101100000", "0101000100000000", "0101011001000000", "0101011110010000", "0101010111100000", "0101010110000000", "0101100010100000", "0101100000100000", "0101101001110000", "0101100011101000", "0101100100101000", "0101011010100000", "0101101000000000", "0101101101010000", "0101101100001000", "0101101010011000", "0101100011101000", "0101100111111000", "0101101011000000", "0101101100101000", "0101101010001000", "0101101101010000", "0101101010010000", "0101101011011000", "0101101010111000", "0101101000100000", "0101100111110000", "0101100011011000", "0101001001000000", "0101100111100000", "0101100111111000", "0101101001100000", "0101101010010000", "0101101010100000", "0101101010000000", "0101101001111000", "0101101010011000", "0101101001111000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101100111111000", "0101100111111000", "0101101101100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001101000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101011001000", "0101100100100000", "0101000110100000", "0101010110000000", "0101011101010000", "0101011111100000", "0101011110010000", "0101100011000000", "0101100111111000", "0101101001110000", "0101100110110000", "0101100010001000", "0101011100110000", "0101101000100000", "0101101100011000", "0101101011010000", "0101101011011000", "0101100010011000", "0101011111110000", "0101100100001000", "0101100110111000", "0101101001010000", "0101101100010000", "0101101100110000", "0101101100001000", "0101101011001000", "0101101001000000", "0101100110100000", "0101100101010000", "0101010010010000", "0101100111101000", "0101101001011000", "0101101011001000", "0101101010010000", "0101101010100000", "0101101011010000", "0101101010000000", "0101101001101000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101000000000", "0101100111111000", "0101101101100000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001101000", "0101101001011000", "0101101001010000", "0101101001101000", "0101101001111000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101010111000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011011000", "0101101010100000", "0101101001010000", "0101000111100000", "0101010111010000", "0101011110010000", "0101100010100000", "0101100011010000", "0101100001011000", "0101100010101000", "0101100110101000", "0101100101110000", "0101100011101000", "0101011100110000", "0101101000100000", "0101101100111000", "0101101011011000", "0101101100010000", "0101101100101000", "0101101010001000", "0101101001010000", "0101101011001000", "0101101100110000", "0101101100011000", "0101101100100000", "0101101100010000", "0101101011100000", "0101101001011000", "0101100101111000", "0101100100110000", "0101001101000000", "0101100111010000", "0101101011010000", "0101101011101000", "0101101010110000", "0101101010101000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001110000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000000000", "0101101101100000", "0101101001101000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001111000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001110000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011100000", "0101101010111000", "0101010010000000", "0101010111000000", "0101011110010000", "0101100010110000", "0101100010100000", "0101100011110000", "0101100101100000", "0101100111011000", "0101101000101000", "0101100010101000", "0101011100110000", "0101100110111000", "0101101100110000", "0101101011011000", "0101101100010000", "0101101110001000", "0101101101010000", "0101101100000000", "0101101100110000", "0101101101100000", "0101101101000000", "0101101100001000", "0101101010011000", "0101101001100000", "0101101000001000", "0101100110010000", "0101100101001000", "0101010100000000", "0101101000101000", "0101101100100000", "0101101000101000", "0101101010110000", "0101101010011000", "0101101010101000", "0101101010010000", "0101101010101000", "0101101010011000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001100000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101001000000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000110000", "0101101000100000", "0101101000100000", "0101101000101000", "0101101000101000", "0101101000001000", "0101101000001000", "0101101000000000", "0101101101100000", "0101101001110000", "0101101001110000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101001111000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011011000", "0101011101110000", "0101010110110000", "0101011100010000", "0101100010001000", "0101100101011000", "0101100100011000", "0101100111100000", "0101101010000000", "0101101000001000", "0101100001100000", "0101011100000000", "0101101000010000", "0101101101100000", "0101101011001000", "0101101011101000", "0101101100101000", "0101101100010000", "0101101100101000", "0101101100111000", "0101101101011000", "0101101100010000", "0101101100001000", "0101101001010000", "0101101001110000", "0101101000111000", "0101100101100000", "0101100001111000", "0101100110101000", "0101101010001000", "0101101100111000", "0101101010100000", "0101101010101000", "0101101010100000", "0101101010111000", "0101101010011000", "0101101010010000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001010000", "0101101001010000", "0101101001001000", "0101101001001000", "0101101000110000", "0101101000110000", "0101101000110000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000010000", "0101101000010000", "0101101000001000", "0101101101100000", "0101101001110000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010010000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011001000", "0101101010101000", "0101101011010000", "0101100110000000", "0101010111010000", "0101011100010000", "0101100000100000", "0101100100111000", "0101100110111000", "0101101000100000", "0101101000011000", "0101100110011000", "0101100000000000", "0101011101010000", "0101100111100000", "0101101101100000", "0101101011000000", "0101101100001000", "0101101101010000", "0101101100000000", "0101101100110000", "0101101100111000", "0101101100011000", "0101101101001000", "0101101100000000", "0101101001111000", "0101101001011000", "0101101001111000", "0101100110100000", "0101100001100000", "0101101001001000", "0101101010111000", "0101100111100000", "0101101010011000", "0101101010111000", "0101101011001000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010101000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000111000", "0101101000100000", "0101101000011000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000011000", "0101101000001000", "0101101101100000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010101000", "0101101010111000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101011011000", "0101101011000000", "0101101011010000", "0101101010100000", "0101010111010000", "0101011110010000", "0101100001001000", "0101100101000000", "0101100110011000", "0101101000110000", "0101100111101000", "0101100101100000", "0101011100010000", "0101011100000000", "0101101000111000", "0101101101110000", "0101101010100000", "0101101001111000", "0101101010110000", "0101101011101000", "0101101011010000", "0101101100011000", "0101101101101000", "0101101100101000", "0101101100100000", "0101101010100000", "0101101010001000", "0101101001000000", "0101100110110000", "0101100011101000", "0101101001000000", "0101101000010000", "0101100111110000", "0101101011010000", "0101101011000000", "0101101010110000", "0101101010100000", "0101101010110000", "0101101010100000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001011000", "0101101001001000", "0101101001000000", "0101101000111000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000010000", "0101101000000000", "0101101101100000", "0101101001111000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101010001000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101011001000", "0101101010111000", "0101101010110000", "0101010100110000", "0101011011100000", "0101100001101000", "0101100101101000", "0101100111101000", "0101100111111000", "0101100111100000", "0101100100110000", "0101011001100000", "0101011110110000", "0101101001011000", "0101101101111000", "0101101010101000", "0101101100011000", "0101101010011000", "0101101000111000", "0101101010011000", "0101101011001000", "0101101100100000", "0101101101010000", "0101101100100000", "0101101011010000", "0101101001000000", "0101101001001000", "0101100111001000", "0101100110010000", "0101101101001000", "0101101011000000", "0101101010000000", "0101101010110000", "0101101010011000", "0101101010101000", "0101101010111000", "0101101010111000", "0101101010101000", "0101101010111000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001001000", "0101101001001000", "0101101001000000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000000000", "0101101101100000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101010000000", "0101101010001000", "0101101010011000", "0101101010101000", "0101101010111000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101011001000", "0101101011011000", "0101101011001000", "0101101011001000", "0101011010110000", "0101011011000000", "0101100001111000", "0101100101100000", "0101100111110000", "0101101000000000", "0101100111101000", "0101100100000000", "0101011100010000", "0101011010100000", "0101100101100000", "0101101010001000", "0101100111000000", "0101101011001000", "0101101010110000", "0101101010000000", "0101100110101000", "0101101010011000", "0101101011001000", "0101101100110000", "0101101100011000", "0101101010111000", "0101101001101000", "0101101000011000", "0101101000100000", "0101100101011000", "0101101100010000", "0101101101100000", "0101101010101000", "0101101010101000", "0101101011001000", "0101101011000000", "0101101010101000", "0101101010011000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001100000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101000000000", "0101101101011000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001111000", "0101101010001000", "0101101010010000", "0101101010100000", "0101101010110000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101011000000", "0101101011011000", "0101100001110000", "0101011010110000", "0101100001001000", "0101100100011000", "0101100100111000", "0101100111110000", "0101100110110000", "0101100100000000", "0101010111100000", "0100100010000000", "0101011110010000", "0101100111111000", "0101011010110000", "0101010000000000", "0101100110111000", "0101101011011000", "0101101000100000", "0101100111001000", "0101101001100000", "0101101011010000", "0101101010100000", "0101101001101000", "0101101001001000", "0101101001110000", "0101100111110000", "0101100111110000", "0101101100011000", "0101101100010000", "0101101010111000", "0101101011000000", "0101101010101000", "0101101010100000", "0101101010101000", "0101101011010000", "0101101011001000", "0101101010100000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001101000", "0101101001101000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000010000", "0101101000010000", "0101101000000000", "0101101101011000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101010001000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010111000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011010000", "0101101010111000", "0101100011000000", "0101010110110000", "0101011110100000", "0101100011011000", "0101100101011000", "0101100111110000", "0101100100100000", "0101100011100000", "0101010100110000", "0101001110000000", "0101011101010000", "0101011110100000", "0101100101000000", "0101100110000000", "0101101010100000", "0101101011110000", "0101101011011000", "0101100011000000", "0101101000101000", "0101101001011000", "0101101001110000", "0101101000101000", "0101100110000000", "0101101001010000", "0101100111110000", "0101100111100000", "0101101101101000", "0101100111001000", "0101101010101000", "0101101011001000", "0101101010011000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001110000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101000110000", "0101101000101000", "0101101000101000", "0101101000100000", "0101101000100000", "0101101000100000", "0101101000001000", "0101101101100000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010100000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011010000", "0101101010101000", "0101101011011000", "0101101011100000", "0101100010011000", "0101010110110000", "0101011010010000", "0101100001011000", "0101100100001000", "0101100101111000", "0101100100111000", "0101100001111000", "0101011101110000", "0101011010100000", "0101010111000000", "0101100011100000", "0101101000001000", "0101101100111000", "0101101100010000", "0101101011101000", "0101101011100000", "0101101000101000", "0101100011111000", "0101100111000000", "0101100111011000", "0101100111100000", "0101100110100000", "0101101000110000", "0101100111111000", "0101100110111000", "0101100110010000", "0101101010110000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001100000", "0101101001100000", "0101101001010000", "0101101000110000", "0101101000100000", "0101101000101000", "0101101000100000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101101100000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011011000", "0101101011100000", "0101101011011000", "0101101011011000", "0101100011001000", "0101011000000000", "0101010110000000", "0101011101000000", "0101100011010000", "0101100101001000", "0101100011101000", "0101100010000000", "0101100011000000", "0101100001011000", "0101100011001000", "0101101001000000", "0101101001101000", "0101101011010000", "0101101100101000", "0101101011111000", "0101101011100000", "0101101010010000", "0101101000010000", "0101100011010000", "0101100110100000", "0101101000010000", "0101101001111000", "0101101001001000", "0101100111101000", "0101100101001000", "0101101010101000", "0101101011101000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001010000", "0101101000111000", "0101101000101000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101101100000", "0101101010010000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101010110000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011110000", "0101101011001000", "0101100111100000", "0101010111010000", "0101010111100000", "0101010111010000", "0101100000110000", "0101100011101000", "0101100001001000", "0101100010000000", "0101100010110000", "0101100100010000", "0101101001001000", "0101101011101000", "0101101011001000", "0101101101001000", "0101101101110000", "0101101101010000", "0101101100100000", "0101101100001000", "0101101010100000", "0101101010010000", "0101101001101000", "0101101010110000", "0101101001100000", "0101101001011000", "0101100111100000", "0101100011011000", "0101101011100000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001011000", "0101101001000000", "0101101000110000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101000010000", "0101101000010000", "0101101101100000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101010110000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011111000", "0101101011000000", "0101101011011000", "0101101011100000", "0101101010111000", "0101010110100000", "0101011000110000", "0101011010100000", "0101100000111000", "0101100010010000", "0101011110010000", "0101011111010000", "0101100011000000", "0101100101000000", "0101101000000000", "0101101010110000", "0101101011100000", "0101101011111000", "0101101100101000", "0101101100010000", "0101101010111000", "0101101001111000", "0101101011100000", "0101101011110000", "0101101100110000", "0101101011101000", "0101101010000000", "0101101000110000", "0101100111000000", "0101100011111000", "0101101010111000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101000100000", "0101101000100000", "0101101000010000", "0101101000010000", "0101101101100000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101010111000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101010101000", "0101101011101000", "0101101011010000", "0101101011010000", "0101101011110000", "0101010111000000", "0101011001110000", "0101011100110000", "0101100011010000", "0101100001100000", "0101010110100000", "0101011010110000", "0101011000110000", "0101010100010000", "0101010100010000", "0101011000010000", "0101011101000000", "0101011001010000", "0101010001000000", "0101010110110000", "0101100000100000", "0101100001100000", "0101100110100000", "0101101011100000", "0101101101000000", "0101101010100000", "0101101010110000", "0101101000001000", "0101100111001000", "0101100001100000", "0101101011010000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010000000", "0101101001110000", "0101101001110000", "0101101001110000", "0101101001011000", "0101101001010000", "0101101001001000", "0101101000110000", "0101101000101000", "0101101000011000", "0101101000011000", "0101101101101000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010110000", "0101101010111000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011110000", "0101101011010000", "0101101011001000", "0101101011110000", "0101101011011000", "0101010110100000", "0101011001110000", "0101011010010000", "0101100101010000", "0101100011011000", "0101010110100000", "0100111000000000", "0100100010000000", "0101100000011000", "0101100101001000", "0101100111001000", "0101101001110000", "0101100110110000", "0101100001110000", "0101100010100000", "0101100100101000", "0101101010100000", "0101100011111000", "0101101010111000", "0101101100111000", "0101101010001000", "0101101001111000", "0101100110000000", "0101100110111000", "0101100001100000", "0101101010111000", "0101101011010000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001100000", "0101101001100000", "0101101001010000", "0101101000111000", "0101101000110000", "0101101000100000", "0101101000011000", "0101101101101000", "0101101010011000", "0101101010011000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011001000", "0101101011010000", "0101101011110000", "0101101011011000", "0101101011100000", "0101010001100000", "0101011001110000", "0101011001110000", "0101100011100000", "0101100111011000", "0101100011001000", "0101010110000000", "0101010011100000", "0101011111010000", "0101011010100000", "0101011000000000", "0101100010100000", "0101100111101000", "0101101001010000", "0101100101101000", "0101101010110000", "0101101101111000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101010010000", "0101101001000000", "0101100100001000", "0101100100101000", "0101100101111000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001000000", "0101101000111000", "0101101000101000", "0101101000100000", "0101101101101000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010110000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011111000", "0101101011100000", "0101101011110000", "0101101011100000", "0101101001011000", "0101010110100000", "0101011010100000", "0101011110110000", "0101101000110000", "0101100011100000", "0101011000100000", "0101010101000000", "0101011111110000", "0101100011000000", "0101100100010000", "0101100111010000", "0101101001010000", "0101101000010000", "0101101001000000", "0101101101110000", "0101101110000000", "0101101101100000", "0101101010110000", "0101101001001000", "0101101010101000", "0101100110111000", "0101100110000000", "0101100011000000", "0101100101011000", "0101101101000000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010011000", "0101101010000000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001000000", "0101101001000000", "0101101000101000", "0101101000100000", "0101101101101000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010100000", "0101101010101000", "0101101010110000", "0101101011000000", "0101101011001000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011101000", "0101101011111000", "0101101011100000", "0101101100001000", "0101101011110000", "0101101011101000", "0101101011111000", "0101101011101000", "0101010110010000", "0101011000010000", "0101010111110000", "0101100011101000", "0101100100000000", "0101100000001000", "0101010110110000", "0101011110100000", "0101011110110000", "0101100011000000", "0101100011101000", "0101100101001000", "0101101001011000", "0101101100111000", "0101101101000000", "0101101101001000", "0101101011100000", "0101101010000000", "0101100111100000", "0101101001001000", "0101100101010000", "0101100100000000", "0101011110010000", "0101100110100000", "0101100001110000", "0101010010110000", "0101101011011000", "0101101011101000", "0101101011111000", "0101101011000000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010000000", "0101101001101000", "0101101001011000", "0101101001011000", "0101101001011000", "0101101001000000", "0101101000110000", "0101101000101000", "0101101101011000", "0101101010011000", "0101101010100000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011110000", "0101101011101000", "0101101011110000", "0101101100000000", "0101101100010000", "0101101100000000", "0101101100010000", "0101101011110000", "0101101100001000", "0101101011111000", "0101010101100000", "0101010110000000", "0101010101000000", "0101011110010000", "0101100011110000", "0101100000111000", "0101011010110000", "0101011010100000", "0101100010101000", "0101100000000000", "0101100010110000", "0101100100010000", "0101101100001000", "0101101100010000", "0101101101101000", "0101101011110000", "0101101011101000", "0101101001011000", "0101101000010000", "0101101000101000", "0101100101001000", "0101100011100000", "0101100101101000", "0101100110100000", "0101010111100000", "0101101111010000", "0101100001010000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101100000000", "0101101010111000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010010000", "0101101010000000", "0101101001110000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101101100000", "0101101010011000", "0101101010101000", "0101101010110000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100001000", "0101101100000000", "0101101011100000", "0101101100001000", "0101101100011000", "0101101011100000", "0101101100011000", "0101101100010000", "0101010101110000", "0101011011010000", "0101010110100000", "0101100000101000", "0101100001100000", "0101100001101000", "0101100000101000", "0101100011111000", "0101100100110000", "0101100111111000", "0101101011101000", "0101101101001000", "0101101101100000", "0101101100101000", "0101101100000000", "0101101011101000", "0101101010110000", "0101101010011000", "0101100111000000", "0101100010111000", "0101100000101000", "0101101000101000", "0101101000000000", "0101011101010000", "0101101111111000", "0101000100100000", "0101101010111000", "0101101011010000", "0101101100000000", "0101101011011000", "0101101011101000", "0101101011111000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101010001000", "0101101010001000", "0101101010000000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001000000", "0101101000111000", "0101101101011000", "0101101010100000", "0101101010110000", "0101101010111000", "0101101011000000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011100000", "0101101011101000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100001000", "0101101100001000", "0101101100010000", "0101101100010000", "0101101100010000", "0101101100010000", "0101101100011000", "0101101100000000", "0101101100100000", "0101101100011000", "0101101100000000", "0101101100110000", "0101101001011000", "0101010110010000", "0101010111110000", "0101011111000000", "0101100001110000", "0101100010001000", "0101100100000000", "0101100110111000", "0101101000101000", "0101101010101000", "0101101011100000", "0101101100111000", "0101101101001000", "0101101100011000", "0101101100110000", "0101101011010000", "0101101000011000", "0101101001000000", "0101100101110000", "0101011100100000", "0101101000001000", "0101101001011000", "0101101010000000", "0101100011001000", "0101101111110000", "0101000010000000", "0101001000000000", "0101101100000000", "0101101011100000", "0101101011011000", "0101101011101000", "0101101011111000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001011000", "0101101001000000", "0101101000111000", "0101101101011000", "0101101010110000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011001000", "0101101011001000", "0101101011011000", "0101101011101000", "0101101011110000", "0101101100001000", "0101101100001000", "0101101100010000", "0101101100010000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100010000", "0101101100010000", "0101101100010000", "0101101101000000", "0101101011101000", "0101101100100000", "0101101100100000", "0101101100000000", "0101101100011000", "0101010010110000", "0101011000100000", "0101011010110000", "0101100010000000", "0101100011111000", "0101100100101000", "0101100101110000", "0101101001100000", "0101101001111000", "0101101100011000", "0101101101110000", "0101101101000000", "0101101101000000", "0101101001110000", "0101101001000000", "0101100110011000", "0101100101000000", "0101100011010000", "0101100110001000", "0101101000100000", "0101101001010000", "0101101001100000", "0101100010101000", "0101101111110000", "0101000011100000", "0100111101000000", "0101101100100000", "0101101011111000", "0101101100010000", "0101101011110000", "0101101011000000", "0101101011110000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101101100000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011010000", "0101101011100000", "0101101011110000", "0101101011111000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100101000", "0101101100000000", "0101101100101000", "0101101100110000", "0101101100011000", "0101101100100000", "0101101100000000", "0101101101011000", "0101000011100000", "0101010110000000", "0101010100010000", "0101100000001000", "0101100010101000", "0101100101111000", "0101100111001000", "0101101000110000", "0101101001000000", "0101101000111000", "0101101100001000", "0101100111101000", "0101101011111000", "0101101000110000", "0101100100000000", "0101100100110000", "0101100010110000", "0101100010001000", "0101101000010000", "0101101011000000", "0101101010110000", "0101101010110000", "0101011101010000", "0101101111101000", "0100111110000000", "0101000100100000", "0100110010000000", "0101101011110000", "0101101011001000", "0101101011110000", "0101101011110000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011011000", "0101101011001000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001100000", "0101101001000000", "0101101000111000", "0101101000110000", "0101101101011000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011101000", "0101101011110000", "0101101011111000", "0101101100001000", "0101101100011000", "0101101100100000", "0101101100011000", "0101101100011000", "0101101100100000", "0101101100100000", "0101101100100000", "0101101100010000", "0101101100011000", "0101101100110000", "0101101100100000", "0101101100010000", "0101101100110000", "0101101101001000", "0100100000000000", "0101100000110000", "0101010001100000", "0101010101010000", "0101010111100000", "0101100000010000", "0101100001110000", "0101100101100000", "0101100110101000", "0101100111101000", "0101101000110000", "0101101000011000", "0101101000101000", "0101101000101000", "0101100101111000", "0101100011010000", "0101100001111000", "0101100010101000", "0101101000010000", "0101101001011000", "0101101001111000", "0101101011001000", "0101100111011000", "0101101111101000", "0101101111111000", "0101000010000000", "0101000110100000", "0100101010000000", "0100011000000000", "0101101100101000", "0101101011011000", "0101101011110000", "0101101011011000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010110000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001001000", "0101101000111000", "0101101000110000", "0101101101011000", "0101101010111000", "0101101011000000", "0101101011010000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011110000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100011000", "0101101100100000", "0101101100100000", "0101101100100000", "0101101100101000", "0101101100101000", "0101101100101000", "0101101100110000", "0101101100101000", "0101101100010000", "0101101100110000", "0101101100101000", "0101101100100000", "0011110000000000", "0100010100000000", "0101100010100000", "0101010100100000", "0101010001110000", "0101011000000000", "0101010110010000", "0101100001101000", "0101100010101000", "0101100101100000", "0101101000101000", "0101100101110000", "0101101000110000", "0101100100110000", "0101100100111000", "0101100100001000", "0101100000111000", "0101100010010000", "0101100111110000", "0101101010001000", "0101101010101000", "0101101011010000", "0101101010100000", "0101100101010000", "0101101111111000", "0101101111101000", "0101000011000000", "0101000110000000", "0100111100000000", "0100110001000000", "0100101100000000", "0101101011110000", "0101101011110000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011010000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001001000", "0101101000111000", "0101101101100000", "0101101010111000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101010110000", "0101101011110000", "0101101100001000", "0101101100000000", "0101101100001000", "0101101100011000", "0101101100001000", "0101101100100000", "0101101100010000", "0101101100011000", "0101101100101000", "0101101100100000", "0101101100111000", "0101101100101000", "0101101100100000", "0101101100101000", "0101101101010000", "0101010010100000", "0100000000000000", "0100110000000000", "0100010000000000", "0101100011100000", "0101011101100000", "0101000100000000", "0101010010110000", "0101011010000000", "0101011010000000", "0101011101000000", "0101100010101000", "0101100010010000", "0101100011110000", "0101100000110000", "0101011111100000", "0101011111110000", "0101100001110000", "0101100010011000", "0101101000000000", "0101101010011000", "0101101011001000", "0101101011111000", "0101101010000000", "0101101000010000", "0101101110011000", "0101101111111000", "0101101111100000", "0101000101100000", "0101001001000000", "0100111111000000", "0100111000000000", "0100111010000000", "0100100110000000", "0101101011001000", "0101101100001000", "0101101011101000", "0101101011100000", "0101101011010000", "0101101011011000", "0101101011110000", "0101101011011000", "0101101010111000", "0101101011011000", "0101101011010000", "0101101010110000", "0101101011011000", "0101101010110000", "0101101011000000", "0101101011000000", "0101101010101000", "0101101010011000", "0101101010100000", "0101101010011000", "0101101010011000", "0101101010010000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101001101000", "0101101001110000", "0101101001011000", "0101101001000000", "0101101101011000", "0101101011001000", "0101101011001000", "0101101011010000", "0101101011010000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011010000", "0101101100000000", "0101101011101000", "0101101011101000", "0101101100011000", "0101101100100000", "0101101100101000", "0101101100010000", "0101101100100000", "0101101100011000", "0101101101001000", "0101101100010000", "0101101100011000", "0101101100010000", "0101101100100000", "0101101101101000", "0000000000000000", "0100100110000000", "0100100010000000", "0100011000000000", "0100011000000000", "0100100000000000", "0101100101001000", "0101100011110000", "0101000101000000", "0101010001100000", "0101010110100000", "0101011100100000", "0101011000110000", "0101011010000000", "0101011111000000", "0101011100110000", "0101011110110000", "0101011110010000", "0101100000000000", "0101100001111000", "0101100111000000", "0101101010110000", "0101101011111000", "0101101100010000", "0101101011111000", "0101101001000000", "0101100100110000", "0101101111111000", "0101101111110000", "0101101111010000", "0101001000000000", "0101000101000000", "0101000110000000", "0101000001000000", "0101000001000000", "0101000001000000", "0100111111000000", "0100111111000000", "0101100000101000", "0101101100011000", "0101101011110000", "0101101011010000", "0101101010111000", "0101101011000000", "0101101011001000", "0101101011001000", "0101101011011000", "0101101011010000", "0101101011001000", "0101101011010000", "0101101011101000", "0101101010100000", "0101101010001000", "0101101011000000", "0101101010100000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001111000", "0101101001101000", "0101101001101000", "0101101001011000", "0101101001000000", "0101101101100000", "0101101011001000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011000000", "0101101011010000", "0101101011100000", "0101101011011000", "0101101011101000", "0101101100011000", "0101101100001000", "0101101100000000", "0101101011110000", "0101101101001000", "0101101100101000", "0101101100001000", "0101101101000000", "0101101100100000", "0101101100011000", "0101101100111000", "0101100001001000", "0100101010000000", "0100101100000000", "0100100110000000", "0100010100000000", "0100100000000000", "0100100010000000", "0100100100000000", "0101100111010000", "0101100111101000", "0101001011100000", "0101010010010000", "0101010101100000", "0101011000100000", "0101011011100000", "0101011111000000", "0101011111110000", "0101100000100000", "0101100001010000", "0101100000010000", "0101100010100000", "0101100110111000", "0101101000110000", "0101101011000000", "0101101011110000", "0101101100101000", "0101101010110000", "0101100111011000", "0101101111001000", "0101101111111000", "0101101111100000", "0101101110111000", "0101000100100000", "0101001011100000", "0101000100000000", "0101000101000000", "0101000001100000", "0101000100000000", "0100111110000000", "0101000111100000", "0101000101100000", "0101000101100000", "0100111001000000", "0101101011101000", "0101101011100000", "0101101011010000", "0101101011011000", "0101101011110000", "0101101011010000", "0101101011011000", "0101101011000000", "0101101011000000", "0101101010101000", "0101101011010000", "0101101011011000", "0101101010011000", "0101101010100000", "0101101010010000", "0101101010010000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001010000", "0101101001000000", "0101101101100000", "0101101011001000", "0101101011010000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011011000", "0101101011010000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011111000", "0101101011100000", "0101101100000000", "0101101011111000", "0101101100100000", "0101101100101000", "0101101100111000", "0101101100011000", "0101101100101000", "0101101100111000", "0101101100001000", "0101101100101000", "0101100111010000", "0100011100000000", "0100101000000000", "0100101000000000", "0100100000000000", "0100010000000000", "0100011000000000", "0100100000000000", "0100010100000000", "0100100010000000", "0101101000011000", "0101101010000000", "0101100101001000", "0101010101010000", "0101011000010000", "0101011010110000", "0101011100010000", "0101011111000000", "0101100000100000", "0101100000100000", "0101100000001000", "0101100011001000", "0101100111000000", "0101101000010000", "0101101001110000", "0101101011010000", "0101101101001000", "0101101011100000", "0101101000000000", "0101100100011000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101110110000", "0101001001100000", "0101000111000000", "0101000101100000", "0101000101000000", "0101000101000000", "0101000101100000", "0101000000100000", "0101000111000000", "0101000111100000", "0101001001000000", "0101001000100000", "0101000111100000", "0101000000000000", "0101100101011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011100000", "0101101011000000", "0101101011010000", "0101101010101000", "0101101010110000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001101000", "0101101001100000", "0101101001010000", "0101101001001000", "0101101001000000", "0101101101100000", "0101101011001000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011010000", "0101101011110000", "0101101011001000", "0101101011110000", "0101101100010000", "0101101100001000", "0101101101001000", "0101101100001000", "0101101100101000", "0101101100101000", "0101101100100000", "0101101100101000", "0101101010011000", "0100100010000000", "0100101010000000", "0100101100000000", "0100110011000000", "0100100010000000", "0100101010000000", "0100100110000000", "0100011100000000", "0100010000000000", "0100100110000000", "0100100000000000", "0101101000110000", "0101101100100000", "0101101010100000", "0101010111010000", "0101011111110000", "0101011111010000", "0101100000010000", "0101100000001000", "0101100001010000", "0101100011010000", "0101100011101000", "0101100101000000", "0101101000010000", "0101101010001000", "0101101010000000", "0101101011100000", "0101101011100000", "0101101010001000", "0101100110010000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101110100000", "0101000111100000", "0101000110100000", "0101000110100000", "0101000110100000", "0101000111000000", "0101000111100000", "0101000000100000", "0101000111000000", "0101000111000000", "0101000101000000", "0101001000000000", "0101000110000000", "0101001000000000", "0101000111000000", "0101000101100000", "0101100110101000", "0101101011001000", "0101101011100000", "0101101011001000", "0101101011101000", "0101101010111000", "0101101011001000", "0101101011000000", "0101101010111000", "0101101010111000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101001111000", "0101101001110000", "0101101001110000", "0101101001100000", "0101101001010000", "0101101001000000", "0101101000111000", "0101101101100000", "0101101011010000", "0101101011011000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101100010000", "0101101011101000", "0101101011101000", "0101101011111000", "0101101100011000", "0101101011111000", "0101101100111000", "0101101100010000", "0101101101000000", "0101101100111000", "0000000000000000", "0100101000000000", "0100101100000000", "0100110000000000", "0100101000000000", "0100100100000000", "0100101110000000", "0100010000000000", "0100011100000000", "0100001000000000", "0100100000000000", "0100101000000000", "0100011000000000", "0101101001101000", "0101101100011000", "0101101101001000", "0101011100100000", "0101100000110000", "0101100010110000", "0101100001001000", "0101100010100000", "0101100001111000", "0101100100100000", "0101100101100000", "0101100111111000", "0101101000101000", "0101101001101000", "0101101011011000", "0101101011011000", "0101101010011000", "0101101000001000", "0101100110111000", "0101101111011000", "0101101111111000", "0101101111111000", "0101101111010000", "0101101110111000", "0101000111100000", "0101000111000000", "0101000110000000", "0101000101100000", "0101000100000000", "0101000111100000", "0101000000100000", "0101000010000000", "0101000110000000", "0101001000000000", "0101000100100000", "0101001000100000", "0101001000000000", "0101000100100000", "0101001010000000", "0101001000100000", "0100111001000000", "0101101100000000", "0101101011101000", "0101101011011000", "0101101011011000", "0101101011001000", "0101101011010000", "0101101010111000", "0101101010111000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010000000", "0101101010000000", "0101101001111000", "0101101001101000", "0101101001011000", "0101101001001000", "0101101001000000", "0101101101100000", "0101101011010000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011110000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011010000", "0101101011000000", "0101101011111000", "0101101100001000", "0101101100011000", "0101101100100000", "0101101101000000", "0101101100010000", "0101101101000000", "0101100000011000", "0100110001000000", "0100101110000000", "0100110000000000", "0100110000000000", "0100101010000000", "0100101110000000", "0100110001000000", "0100100100000000", "0100101000000000", "0100010100000000", "0100010000000000", "0100011100000000", "0100101100000000", "0100011100000000", "0101101010111000", "0101101101100000", "0101101111000000", "0101101110101000", "0101100001110000", "0101100100001000", "0101100100111000", "0101100011101000", "0101100011010000", "0101100100101000", "0101100111011000", "0101100111000000", "0101101001110000", "0101101001011000", "0101101001100000", "0101101010101000", "0101101000011000", "0101100101100000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101000100000", "0101000111000000", "0101000111000000", "0101000110100000", "0101001000000000", "0101000111000000", "0101000101100000", "0101000010100000", "0100110101000000", "0101000110100000", "0101000111100000", "0101000101100000", "0101000110100000", "0101000110100000", "0101000111100000", "0101000101000000", "0101000111000000", "0101000101100000", "0101000110000000", "0101100010101000", "0101101011101000", "0101101011010000", "0101101011001000", "0101101011001000", "0101101010110000", "0101101010111000", "0101101010100000", "0101101010011000", "0101101010010000", "0101101010001000", "0101101010000000", "0101101010000000", "0101101001110000", "0101101001011000", "0101101001001000", "0101101000111000", "0101101101100000", "0101101011011000", "0101101011101000", "0101101011110000", "0101101011110000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011110000", "0101101011110000", "0101101011110000", "0101101011110000", "0101101011101000", "0101101100000000", "0101101011011000", "0101101011111000", "0101101100010000", "0101101100011000", "0101101100010000", "0101101101010000", "0101011110000000", "0100101110000000", "0100110000000000", "0100110000000000", "0100101110000000", "0100101110000000", "0100110001000000", "0100101100000000", "0100110010000000", "0100101110000000", "0100101010000000", "0100101010000000", "0100010100000000", "0100100000000000", "0100100010000000", "0100110001000000", "0100010100000000", "0101101011100000", "0101101010011000", "0101100101101000", "0101101010101000", "0101101010111000", "0101101100001000", "0101100111000000", "0101100101101000", "0101100101010000", "0101100101000000", "0101100111000000", "0101100111100000", "0101101000001000", "0101101000110000", "0101101000001000", "0101101001000000", "0101100101110000", "0101101111100000", "0101101111100000", "0101101111111000", "0101101111101000", "0101101111110000", "0101101111101000", "0101011110100000", "0101001000100000", "0101000111100000", "0101000111000000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000011000000", "0101000001000000", "0101000101100000", "0101000110000000", "0101000101100000", "0101000101100000", "0101000100100000", "0101000110000000", "0101000111000000", "0101000110000000", "0101000111000000", "0101000111100000", "0101000111000000", "0101000010000000", "0101101100000000", "0101101011100000", "0101101011011000", "0101101011001000", "0101101011000000", "0101101010101000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101010000000", "0101101001111000", "0101101001101000", "0101101001100000", "0101101001001000", "0101101000111000", "0101101101011000", "0101101011100000", "0101101011101000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011011000", "0101101011110000", "0101101011110000", "0101101011100000", "0101101100001000", "0101101011101000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100001000", "0101101100010000", "0101101100101000", "0101101000000000", "0100110001000000", "0100110001000000", "0100101100000000", "0100110000000000", "0100110001000000", "0100110001000000", "0100110010000000", "0100110011000000", "0100110011000000", "0100110001000000", "0100101110000000", "0100011000000000", "0100101100000000", "0100010100000000", "0100100000000000", "0100100100000000", "0100110011000000", "0100010100000000", "0101101111011000", "0101100100100000", "0101100110111000", "0101101010111000", "0101101101011000", "0101101011110000", "0101101010101000", "0101100111110000", "0101100111000000", "0101100101111000", "0101100110000000", "0101100110011000", "0101100110101000", "0101100110001000", "0101100111001000", "0101100110111000", "0101101111101000", "0101101101110000", "0101101100100000", "0101101111100000", "0101101111101000", "0101101111111000", "0101101111111000", "0101010011000000", "0101001010000000", "0101001001000000", "0101001000100000", "0101000111100000", "0101000111100000", "0101000111100000", "0101000011100000", "0101000001000000", "0101000110000000", "0101000110100000", "0101000110000000", "0101000110100000", "0101000110000000", "0101000101100000", "0101000111000000", "0101000111100000", "0101000110100000", "0101001001100000", "0101000111100000", "0101000111000000", "0101001001000000", "0101101010100000", "0101101011011000", "0101101011011000", "0101101010111000", "0101101010111000", "0101101010110000", "0101101010101000", "0101101010001000", "0101101010001000", "0101101010010000", "0101101001101000", "0101101001100000", "0101101001011000", "0101101001001000", "0101101101011000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011101000", "0101101011101000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101011100000", "0101101011110000", "0101101011101000", "0101101100001000", "0101101100001000", "0101101101000000", "0100111011000000", "0100110011000000", "0100101110000000", "0100101110000000", "0100110000000000", "0100110010000000", "0100110011000000", "0100110011000000", "0100110011000000", "0100110011000000", "0100110011000000", "0100110010000000", "0100101110000000", "0100101000000000", "0100011100000000", "0100100100000000", "0100101000000000", "0100101010000000", "0100101100000000", "0100101010000000", "0101101010100000", "0101100110111000", "0101101000001000", "0101101000111000", "0101101101000000", "0101101100001000", "0101101011010000", "0101101101000000", "0101101001000000", "0101100111011000", "0101100110110000", "0101100110000000", "0101100101000000", "0101100101100000", "0101101000101000", "0101101111011000", "0101101010111000", "0101101110000000", "0101101100111000", "0101101011010000", "0101101111111000", "0101101111111000", "0101101111100000", "0101001110000000", "0101001001000000", "0101001000100000", "0101001001000000", "0101001000100000", "0101001000100000", "0101001000000000", "0101000101000000", "0101000011100000", "0101000101100000", "0101000111000000", "0101000110100000", "0101000110100000", "0101000110000000", "0101000110000000", "0101001000000000", "0101001000000000", "0101001001100000", "0101001000000000", "0101001001000000", "0101001001000000", "0101001000100000", "0101000111000000", "0101000101100000", "0101101011111000", "0101101011010000", "0101101011010000", "0101101010010000", "0101101010011000", "0101101010101000", "0101101001111000", "0101101010000000", "0101101010001000", "0101101001101000", "0101101001100000", "0101101001001000", "0101101101100000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011101000", "0101101011110000", "0101101011100000", "0101101011010000", "0101101100000000", "0101101100000000", "0101101100010000", "0101101100001000", "0101101100011000", "0101101000010000", "0000000000000000", "0100110010000000", "0100110000000000", "0100110000000000", "0100110000000000", "0100110100000000", "0100110011000000", "0100110100000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110011000000", "0100110011000000", "0100100100000000", "0100110100000000", "0100100100000000", "0100101010000000", "0100100000000000", "0100100110000000", "0100110011000000", "0101010110000000", "0101101011001000", "0101101001010000", "0101101010110000", "0101101010010000", "0101101100000000", "0101101100010000", "0101101011101000", "0101101100000000", "0101101011110000", "0101101010001000", "0101100111111000", "0101100110111000", "0101100110010000", "0101100101001000", "0101101000011000", "0101101111110000", "0101101110111000", "0101101111001000", "0101101101010000", "0101101010100000", "0101101001101000", "0101101111111000", "0101101111110000", "0101000110100000", "0101001001000000", "0101001000100000", "0101001001100000", "0101001001000000", "0101001000000000", "0101000110100000", "0101000100000000", "0101000100000000", "0101000110000000", "0101001000000000", "0101000111100000", "0101000111000000", "0101000110000000", "0101000110000000", "0101001000000000", "0101000111100000", "0101001000100000", "0101001000000000", "0101000111100000", "0101001001000000", "0101001000000000", "0101000111000000", "0101001001100000", "0101000111100000", "0101000101000000", "0101101011001000", "0101101010100000", "0101101010101000", "0101101010000000", "0101101010101000", "0101101001110000", "0101101001111000", "0101101001111000", "0101101001101000", "0101101001010000", "0101101101100000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101010110000", "0101101100001000", "0101101011111000", "0101101011011000", "0101101100000000", "0101101011111000", "0101101100011000", "0100101100000000", "0100110010000000", "0100110010000000", "0100110000000000", "0100110011000000", "0100110101000000", "0100110000000000", "0100110011000000", "0100110101000000", "0100110110000000", "0100111000000000", "0100110111000000", "0100110110000000", "0100110101000000", "0100110100000000", "0100110100000000", "0100100000000000", "0100110011000000", "0100101000000000", "0100101010000000", "0100101000000000", "0100101100000000", "0100110001000000", "0101100010111000", "0101101100010000", "0101101011011000", "0101101100110000", "0101101100000000", "0101101011111000", "0101101100100000", "0101101100111000", "0101101101100000", "0101101100011000", "0101101100001000", "0101101010001000", "0101101000101000", "0101100111101000", "0101100110101000", "0101101100110000", "0101101111111000", "0101101111110000", "0101101111100000", "0101101101001000", "0101101011011000", "0101101010001000", "0101101111000000", "0101101111100000", "0101001011000000", "0101001001100000", "0101001000000000", "0101001000100000", "0101001000100000", "0101000111000000", "0101000101000000", "0101000011100000", "0101000100100000", "0101000110000000", "0101001000100000", "0101001000000000", "0101000111000000", "0101000101100000", "0101000110000000", "0101000111100000", "0101000111100000", "0101000111000000", "0101001001100000", "0101001100000000", "0101000111100000", "0101001000000000", "0101001000000000", "0101001000000000", "0101000111100000", "0101000111000000", "0101000111100000", "0101100011101000", "0101101011001000", "0101101010010000", "0101101010011000", "0101101010001000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001011000", "0101101101100000", "0101101011111000", "0101101011110000", "0101101011110000", "0101101011101000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011011000", "0101101011111000", "0101101011101000", "0101101011000000", "0101101100010000", "0101101100100000", "0101101011101000", "0101100101001000", "0100110100000000", "0100110100000000", "0100110011000000", "0100110000000000", "0100111000000000", "0100110010000000", "0100101100000000", "0100110110000000", "0100110101000000", "0100110101000000", "0100110111000000", "0100111001000000", "0100111000000000", "0100110111000000", "0100110111000000", "0100110110000000", "0100110100000000", "0100101100000000", "0100110000000000", "0100101010000000", "0100101100000000", "0100101110000000", "0100101110000000", "0100110110000000", "0101100100111000", "0101101101000000", "0101101100110000", "0101101101110000", "0101101101011000", "0101101100011000", "0101101100100000", "0101101101000000", "0101101110000000", "0101101100010000", "0101101100100000", "0101101100010000", "0101101010000000", "0101100111101000", "0101100111101000", "0101101101010000", "0101101111110000", "0101101111111000", "0101101111101000", "0101101100111000", "0101101100011000", "0101101010110000", "0101101010010000", "0101101111010000", "0101001000100000", "0101001001000000", "0101000111000000", "0101001000000000", "0101001000000000", "0101000111100000", "0101000110000000", "0101000100000000", "0101000101100000", "0101000101000000", "0101000111100000", "0101000111000000", "0101000110100000", "0101000101100000", "0101000110100000", "0101001000100000", "0101001000000000", "0101001001100000", "0101001000100000", "0101000111100000", "0101000101100000", "0101000111100000", "0101001001100000", "0101001001000000", "0101000111100000", "0101001000000000", "0101000111000000", "0101000111000000", "0101011001100000", "0101101010111000", "0101101010011000", "0101101010101000", "0101101010001000", "0101101001111000", "0101101001110000", "0101101001011000", "0101101101101000", "0101101100000000", "0101101100000000", "0101101011111000", "0101101011110000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011000000", "0101101100001000", "0101101011100000", "0101101011110000", "0101101011101000", "0101101100010000", "0100111110000000", "0100110001000000", "0100110010000000", "0100110101000000", "0100110011000000", "0100110110000000", "0100110010000000", "0100111001000000", "0100110010000000", "0100110101000000", "0100110101000000", "0100111000000000", "0100111001000000", "0100110111000000", "0100110111000000", "0100111001000000", "0100110111000000", "0100110011000000", "0100110101000000", "0100110001000000", "0100101110000000", "0100101110000000", "0100100010000000", "0100100100000000", "0101000010000000", "0101100011011000", "0101101111010000", "0101101110001000", "0101101110111000", "0101101110101000", "0101101100111000", "0101101100100000", "0101101100100000", "0101101011111000", "0101101100101000", "0101101100000000", "0101101011111000", "0101101010000000", "0101101000101000", "0101101000010000", "0101101000110000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101110000000", "0101101110000000", "0101101100110000", "0101101010110000", "0101101111100000", "0101001010000000", "0101001001100000", "0101000111100000", "0101000111100000", "0101001000000000", "0101000111100000", "0101000110000000", "0101000100000000", "0101000100100000", "0101000101100000", "0101000111000000", "0101000110100000", "0101000110100000", "0101000110000000", "0101000110100000", "0101001000100000", "0101001000000000", "0101000111000000", "0101001000100000", "0101001001100000", "0101000111100000", "0101001001000000", "0101000110100000", "0101000101000000", "0101001000000000", "0101001000000000", "0101000110100000", "0101001000000000", "0101001000000000", "0101000100100000", "0101101011010000", "0101101010110000", "0101101010000000", "0101101001111000", "0101101001110000", "0101101001011000", "0101101101101000", "0101101100000000", "0101101011111000", "0101101011110000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101100000000", "0101101011111000", "0101101100001000", "0101101011110000", "0101101100001000", "0101100101011000", "0100111000000000", "0100110100000000", "0100110100000000", "0100110111000000", "0100110111000000", "0100110010000000", "0100110100000000", "0100110010000000", "0100110101000000", "0100111000000000", "0100110101000000", "0100111001000000", "0100111001000000", "0100110110000000", "0100110111000000", "0100111011000000", "0100111000000000", "0100110001000000", "0100111000000000", "0100110000000000", "0100110000000000", "0100101100000000", "0100100110000000", "0100101100000000", "0101000010100000", "0101100000011000", "0101101111011000", "0101101111100000", "0101101111011000", "0101101110111000", "0101101110000000", "0101101100111000", "0101101100110000", "0101101101110000", "0101101100001000", "0101101100000000", "0101101011001000", "0101101001111000", "0101101001011000", "0101101001010000", "0101101000001000", "0101101111011000", "0101101111111000", "0101101111100000", "0101101111001000", "0101101110000000", "0101101101110000", "0101101100010000", "0101101111101000", "0101001000000000", "0101001001100000", "0101001000000000", "0101001000100000", "0101001000000000", "0101000111000000", "0101000101100000", "0101000011000000", "0101000010100000", "0101000111000000", "0101000111100000", "0101000110100000", "0101000110100000", "0101000110100000", "0101000110100000", "0101001000000000", "0101000111100000", "0101001010000000", "0101000110100000", "0101000110100000", "0101000111100000", "0101000111100000", "0101001000000000", "0101001000000000", "0101000111000000", "0101000111100000", "0101000100000000", "0101001000100000", "0101001001100000", "0101000001000000", "0101000010100000", "0101101010010000", "0101101010011000", "0101101010000000", "0101101001111000", "0101101001100000", "0101101101101000", "0101101011110000", "0101101011110000", "0101101011101000", "0101101011100000", "0101101011011000", "0101101011011000", "0101101011101000", "0101101011110000", "0101101011111000", "0101101011110000", "0101101011111000", "0101101011111000", "0101101100001000", "0100100000000000", "0100111110000000", "0100110011000000", "0100111000000000", "0100110010000000", "0100110010000000", "0100111001000000", "0100110100000000", "0100110100000000", "0100110111000000", "0100110101000000", "0100110101000000", "0100111001000000", "0100111000000000", "0100110101000000", "0100110111000000", "0100111100000000", "0100111000000000", "0100110000000000", "0100110110000000", "0100110001000000", "0100110101000000", "0100101000000000", "0100101100000000", "0100110010000000", "0101000010100000", "0101100001001000", "0101101111101000", "0101101111101000", "0101101111101000", "0101101111101000", "0101101111000000", "0101101100101000", "0101101100000000", "0101101100110000", "0101101011100000", "0101101100011000", "0101101011111000", "0101101010111000", "0101101001000000", "0101101000100000", "0101100110111000", "0101100100011000", "0101101111101000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101110101000", "0101101101000000", "0101101111100000", "0101000100000000", "0101001000000000", "0101000111100000", "0101001000100000", "0101001000100000", "0101000111100000", "0101000110000000", "0101000011000000", "0101000010100000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000111000000", "0101000111100000", "0101000111100000", "0101001000100000", "0101001000100000", "0101001000100000", "0101000111100000", "0101001000000000", "0101000111100000", "0101000110000000", "0101001001100000", "0101000101100000", "0101000111000000", "0101000101100000", "0101000111000000", "0101001001100000", "0101000110000000", "0101000010000000", "0100111111000000", "0101101010101000", "0101101010011000", "0101101010000000", "0101101001111000", "0101101001100000", "0101101101101000", "0101101011110000", "0101101011101000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011110000", "0101101011111000", "0101101100000000", "0101101011110000", "0101101100010000", "0101101011110000", "0101101100011000", "0101101100100000", "0100110010000000", "0101000001000000", "0100110011000000", "0100110100000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110101000000", "0100110111000000", "0100111000000000", "0100110111000000", "0100111000000000", "0100110011000000", "0100111001000000", "0100111000000000", "0100111010000000", "0100111011000000", "0100111001000000", "0100101110000000", "0100110101000000", "0100110010000000", "0100110000000000", "0100101000000000", "0100101010000000", "0100101010000000", "0101000011100000", "0101011010100000", "0101101111110000", "0101101111111000", "0101101111011000", "0101101111111000", "0101101111101000", "0101101101111000", "0101101100010000", "0101101100101000", "0101101100010000", "0101101011100000", "0101101010110000", "0101101010011000", "0101101001111000", "0101101000111000", "0101100110011000", "0101100011010000", "0101101111011000", "0101101111111000", "0101101111110000", "0101101111011000", "0101101111101000", "0101101110100000", "0101101101000000", "0101001000000000", "0101001010000000", "0101000111100000", "0101001000100000", "0101001000100000", "0101000110100000", "0101000100100000", "0101000100000000", "0101000110000000", "0101000111000000", "0101000110000000", "0101000110000000", "0101000101100000", "0101001000000000", "0101001001100000", "0101000110100000", "0101001000000000", "0101000111100000", "0101000111000000", "0101000110100000", "0101000111000000", "0101000111100000", "0101001000000000", "0101000111100000", "0101000111000000", "0101000101100000", "0101000111100000", "0101000100100000", "0101000101100000", "0101000000000000", "0100110101000000", "0101101010111000", "0101101010100000", "0101101010010000", "0101101001111000", "0101101001110000", "0101101101011000", "0101101011100000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011101000", "0101101011110000", "0101101011111000", "0101101100000000", "0101101100010000", "0101101100010000", "0101101100100000", "0101101011101000", "0101101100001000", "0100111000000000", "0100111100000000", "0100110011000000", "0100110100000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110111000000", "0100111000000000", "0100110111000000", "0100110100000000", "0100110100000000", "0100111010000000", "0100111001000000", "0100111100000000", "0100111101000000", "0100111010000000", "0100101000000000", "0100111010000000", "0100101100000000", "0100101110000000", "0100110000000000", "0100100110000000", "0100110111000000", "0101000010100000", "0101011101000000", "0101101111110000", "0101101111111000", "0101101111001000", "0101101111111000", "0101101111111000", "0101101110100000", "0101101100100000", "0101101011101000", "0101101101010000", "0101101100000000", "0101101011100000", "0101101010111000", "0101101001101000", "0101101000110000", "0101100110000000", "0101101011101000", "0101101111001000", "0101101111100000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101110111000", "0101100100011000", "0101000011000000", "0101001001100000", "0101000111000000", "0101001000000000", "0101001000100000", "0101000111100000", "0101000110100000", "0101000101100000", "0101000110100000", "0101000111100000", "0101000111000000", "0101000110000000", "0101000100000000", "0101000110100000", "0101001000100000", "0101000110100000", "0101000111100000", "0101000111100000", "0101000111000000", "0101000110100000", "0101000111000000", "0101000111000000", "0101000110100000", "0101000101000000", "0101000100000000", "0101000101100000", "0101000011000000", "0100101100000000", "0101000100000000", "0100111101000000", "0100110101000000", "0101101010101000", "0101101010010000", "0101101010010000", "0101101010000000", "0101101001110000", "0101101101011000", "0101101011011000", "0101101011011000", "0101101011100000", "0101101011101000", "0101101011110000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101100001000", "0101101011101000", "0101101100100000", "0101101011111000", "0100110111000000", "0100111011000000", "0100110000000000", "0100110100000000", "0100110101000000", "0100110110000000", "0100110101000000", "0100110110000000", "0100110111000000", "0100110111000000", "0100110110000000", "0100110100000000", "0100110111000000", "0100111001000000", "0100110111000000", "0100111011000000", "0100111110000000", "0100111100000000", "0100101010000000", "0100101110000000", "0100111011000000", "0100110000000000", "0100100100000000", "0100101100000000", "0100110010000000", "0101000110000000", "0101101110110000", "0101101111110000", "0101101111110000", "0101101111001000", "0101101111111000", "0101101111111000", "0101101111010000", "0101101101011000", "0101101011100000", "0101101100111000", "0101101011111000", "0101101011100000", "0101101001010000", "0101101010110000", "0101101000110000", "0101100101011000", "0101101110111000", "0101101111111000", "0101101111100000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101010111000000", "0101001001100000", "0101001001100000", "0101000111000000", "0101001000000000", "0101001000100000", "0101001000000000", "0101000111000000", "0101000101100000", "0101000101100000", "0101000110000000", "0101000111000000", "0101000110000000", "0101000100000000", "0101000110000000", "0101001001000000", "0101001000000000", "0101001000000000", "0101000101100000", "0101000100100000", "0101000100100000", "0101000101100000", "0101000110100000", "0101000111000000", "0101000110100000", "0101000110000000", "0101000100100000", "0101000100100000", "0100110010000000", "0101000001100000", "0101000000100000", "0100110010000000", "0101101000101000", "0101101010011000", "0101101010011000", "0101101010000000", "0101101001111000", "0101101101011000", "0101101011100000", "0101101011100000", "0101101011101000", "0101101011110000", "0101101011110000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100000000", "0101101011111000", "0101101100110000", "0101101100010000", "0100110010000000", "0101000010000000", "0100101010000000", "0100110011000000", "0100110101000000", "0100110110000000", "0100110110000000", "0100110110000000", "0100110111000000", "0100110110000000", "0100110101000000", "0100110101000000", "0100111000000000", "0100110111000000", "0100110110000000", "0100111100000000", "0100111111000000", "0100111011000000", "0100110000000000", "0100110101000000", "0100110101000000", "0100101110000000", "0100110000000000", "0100101100000000", "0100110110000000", "0101000101000000", "0101101111100000", "0101101111110000", "0101101111101000", "0101101111011000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101110100000", "0101101100110000", "0101101010011000", "0101101100111000", "0101101100000000", "0101101010101000", "0101101001001000", "0101100111111000", "0101101111100000", "0101101111100000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101000101100000", "0101001001000000", "0101001001000000", "0101000111100000", "0101001000100000", "0101001000100000", "0101000111100000", "0101000111100000", "0101000101100000", "0101000101000000", "0101000101100000", "0101000111000000", "0101000110000000", "0101000101000000", "0101000111000000", "0101001000100000", "0101001000000000", "0101001000000000", "0101000111000000", "0101000101100000", "0101000100000000", "0101000100000000", "0101000101000000", "0101000110000000", "0101000110000000", "0101000110000000", "0101000011000000", "0101000001000000", "0101000010100000", "0101000100000000", "0100110110000000", "0100111001000000", "0101100000101000", "0101101010101000", "0101101010011000", "0101101010001000", "0101101001111000", "0101101101011000", "0101101011110000", "0101101011110000", "0101101011110000", "0101101011110000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100010000", "0101101100010000", "0101101100010000", "0100111000000000", "0100111101000000", "0100100100000000", "0100110011000000", "0100110101000000", "0100110110000000", "0100110101000000", "0100110101000000", "0100110110000000", "0100110110000000", "0100110101000000", "0100110100000000", "0100110110000000", "0100110111000000", "0100111010000000", "0101000000000000", "0101000000100000", "0100110111000000", "0100110010000000", "0100110011000000", "0100110111000000", "0100110011000000", "0100101110000000", "0100101000000000", "0100111001000000", "0101000110100000", "0101101111000000", "0101101111111000", "0101101111101000", "0101101111010000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111010000", "0101101101111000", "0101101100011000", "0101101101110000", "0101101010111000", "0101101010010000", "0101101001101000", "0101101110010000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111010000", "0101000000100000", "0101000110100000", "0101000111100000", "0101000111000000", "0101001000100000", "0101001000000000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000101100000", "0101000111000000", "0101000111100000", "0101000110000000", "0101000110000000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000111000000", "0101001000000000", "0101000110100000", "0101000100000000", "0101000011000000", "0101000011100000", "0101000100100000", "0101000100100000", "0101000101000000", "0101000011000000", "0100111010000000", "0101000100100000", "0100111011000000", "0100111010000000", "0100111000000000", "0101000010100000", "0101101010100000", "0101101010011000", "0101101010001000", "0101101010000000", "0101101101100000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101011111000", "0101101100000000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100001000", "0101101100101000", "0101101011110000", "0101101100100000", "0101101101110000", "0100110111000000", "0100110111000000", "0100101010000000", "0100110010000000", "0100110100000000", "0100110110000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110111000000", "0100111001000000", "0100111111000000", "0101000000100000", "0100110010000000", "0100110111000000", "0100110011000000", "0100110010000000", "0100110010000000", "0100110001000000", "0100101100000000", "0100110101000000", "0101000111000000", "0101101111010000", "0101101111111000", "0101101111101000", "0101101111010000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111011000", "0101101110010000", "0101101101111000", "0101101010011000", "0101101010101000", "0101101010011000", "0101101011110000", "0101101111111000", "0101101111110000", "0101101111100000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111110000", "0101101110111000", "0101001000000000", "0101001001100000", "0101000110100000", "0101000111000000", "0101001000100000", "0101000111000000", "0101000101000000", "0101000110000000", "0101000101100000", "0101000100100000", "0101000111100000", "0101001000000000", "0101000101100000", "0101000110000000", "0101000111100000", "0101000110100000", "0101000110100000", "0101000111100000", "0101000110100000", "0101000101100000", "0101000100000000", "0101000011100000", "0101000100000000", "0101000100100000", "0101000101000000", "0101000101000000", "0101000001100000", "0100101000000000", "0101000001000000", "0100111111000000", "0100111011000000", "0100110011000000", "0100110110000000", "0101101010101000", "0101101010011000", "0101101010001000", "0101101010000000", "0101101101100000", "0101101100000000", "0101101100001000", "0101101100001000", "0101101100010000", "0101101100010000", "0101101100011000", "0101101100011000", "0101101100011000", "0101101100100000", "0101101100011000", "0101101100101000", "0101101100101000", "0101101101101000", "0100101110000000", "0100111101000000", "0100110111000000", "0100110010000000", "0100110100000000", "0100110110000000", "0100110101000000", "0100110100000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110011000000", "0100111000000000", "0100110111000000", "0100111100000000", "0101000000100000", "0100101110000000", "0100111010000000", "0100110011000000", "0100110111000000", "0100110100000000", "0100101010000000", "0100110000000000", "0100111000000000", "0101000101100000", "0101101110111000", "0101101111110000", "0101101111111000", "0101101111100000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111101000", "0101101110111000", "0101101110111000", "0101101100101000", "0101101100111000", "0101101001111000", "0101101111111000", "0101101111011000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101110001000", "0101001001000000", "0101000111100000", "0101000111000000", "0101000111100000", "0101001000100000", "0101000110000000", "0101000100000000", "0101000101100000", "0101000101000000", "0101000100000000", "0101000110100000", "0101001000100000", "0101000101100000", "0101000110000000", "0101000111100000", "0101000111100000", "0101000111100000", "0101000111100000", "0101000110100000", "0101000110000000", "0101000101000000", "0101000100000000", "0101000100000000", "0101000100000000", "0101000100000000", "0101000100000000", "0101000010100000", "0101000001100000", "0101000010000000", "0101000011100000", "0100110110000000", "0100110100000000", "0100110110000000", "0101101010010000", "0101101010011000", "0101101010001000", "0101101010000000", "0101101101100000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100100000", "0101101100100000", "0101101100100000", "0101101100011000", "0101101100010000", "0101101100101000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101000010000", "0100110110000000", "0100110110000000", "0100111101000000", "0100110010000000", "0100110101000000", "0100110110000000", "0100110101000000", "0100110100000000", "0100110101000000", "0100110110000000", "0100110101000000", "0100110010000000", "0100110001000000", "0100111011000000", "0100111000000000", "0100111101000000", "0101000001000000", "0100101000000000", "0100111001000000", "0100110100000000", "0100110110000000", "0100110011000000", "0100101100000000", "0100110000000000", "0100110111000000", "0101000100100000", "0101101111011000", "0101101111100000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101110010000", "0101101100111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111100000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111110000", "0101101111111000", "0101101111100000", "0101101101111000", "0101000111100000", "0101001000100000", "0101000111000000", "0101000111100000", "0101001000100000", "0101000110000000", "0101000100100000", "0101000110100000", "0101000110100000", "0101000101100000", "0101000110000000", "0101001000100000", "0101000110100000", "0101000110000000", "0101000111100000", "0101000111100000", "0101000111000000", "0101000101000000", "0101000110000000", "0101000101000000", "0101000100000000", "0101000011000000", "0101000011000000", "0101000011000000", "0101000011100000", "0101000100000000", "0101000000000000", "0101000000100000", "0101000110100000", "0100111010000000", "0100110110000000", "0100111001000000", "0100110101000000", "0101101010110000", "0101101010011000", "0101101010001000", "0101101010000000", "0101101101100000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100011000", "0101101100100000", "0101101100100000", "0101101100100000", "0101101100100000", "0101101100110000", "0101101100100000", "0101101100110000", "0101101100111000", "0101010101100000", "0100110010000000", "0100111000000000", "0101000001100000", "0100110001000000", "0100110111000000", "0100110110000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110110000000", "0100110101000000", "0100110100000000", "0100110111000000", "0100110111000000", "0100111000000000", "0100111100000000", "0101000001000000", "0100110001000000", "0100111010000000", "0100110101000000", "0100110101000000", "0100110001000000", "0100110001000000", "0100110000000000", "0100111001000000", "0101000100000000", "0101101111011000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111110000", "0101101111110000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101101110000", "0101000101100000", "0101000111000000", "0101000111000000", "0101000111100000", "0101000110000000", "0101000111000000", "0101000101000000", "0101000101100000", "0101000101100000", "0101000101000000", "0101000111000000", "0101000111100000", "0101000110100000", "0101000110000000", "0101000111000000", "0101000111100000", "0101000110000000", "0101000101000000", "0101000100100000", "0101000101100000", "0101000110000000", "0101000100000000", "0101000100100000", "0101000011100000", "0101000011100000", "0101000011000000", "0100110000000000", "0101000001100000", "0101000011000000", "0100111011000000", "0100110011000000", "0100110110000000", "0100111111000000", "0101101010011000", "0101101010100000", "0101101010010000", "0101101010000000", "0101101101100000", "0101101100001000", "0101101100010000", "0101101100011000", "0101101100100000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101100101000", "0101101101101000", "0101101100110000", "0100111010000000", "0100110001000000", "0100111001000000", "0101000011000000", "0100110000000000", "0100110110000000", "0100110101000000", "0100110110000000", "0100110111000000", "0100110111000000", "0100110111000000", "0100110101000000", "0100110011000000", "0100110110000000", "0100110111000000", "0100111010000000", "0100111110000000", "0101000001100000", "0100110011000000", "0100111010000000", "0100110110000000", "0100110100000000", "0100110000000000", "0100110000000000", "0100110000000000", "0100111100000000", "0101000110000000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111010000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111010000", "0101101111110000", "0101101111111000", "0101101111100000", "0101101000101000", "0101000011000000", "0101001010000000", "0101000111100000", "0101000111100000", "0101000110100000", "0101000111100000", "0101000110000000", "0101000110000000", "0101000100000000", "0101000100000000", "0101000111100000", "0101001000100000", "0101000111000000", "0101000110000000", "0101000110100000", "0101000111000000", "0101000110000000", "0101000100100000", "0101000101000000", "0101000101000000", "0101000110000000", "0101000100000000", "0101000100100000", "0101000011100000", "0101000011100000", "0101000001100000", "0100101100000000", "0101000100100000", "0101000000000000", "0100111001000000", "0100110001000000", "0100110110000000", "0100111001000000", "0101101010110000", "0101101010100000", "0101101010010000", "0101101010001000", "0101101101100000", "0101101100010000", "0101101100011000", "0101101100100000", "0101101100101000", "0101101100110000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101101000000", "0101101100111000", "0101101101000000", "0101101100101000", "0100111001000000", "0100110001000000", "0100110010000000", "0101000010000000", "0100101110000000", "0100110100000000", "0100110100000000", "0100110101000000", "0100110111000000", "0100110110000000", "0100110110000000", "0100110100000000", "0100110011000000", "0100110101000000", "0100110110000000", "0100111001000000", "0100111111000000", "0101000010000000", "0100110100000000", "0100111010000000", "0100110111000000", "0100110100000000", "0100110001000000", "0100110000000000", "0100101110000000", "0100111101000000", "0101000101100000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101110000000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111010000", "0101101111111000", "0101101111011000", "0101101111110000", "0101101111011000", "0101010100000000", "0101000111000000", "0101000101100000", "0101001000000000", "0101000111100000", "0101000111100000", "0101000111000000", "0101000111000000", "0101000111000000", "0101000011000000", "0101000101000000", "0101001000000000", "0101001001100000", "0101001000000000", "0101000110000000", "0101000110100000", "0101000111100000", "0101000110000000", "0101000100100000", "0101000101100000", "0101000101000000", "0101000110100000", "0101000101000000", "0101000100000000", "0101000011000000", "0101000011100000", "0101000000100000", "0100111101000000", "0101000011000000", "0101000000100000", "0100111001000000", "0100110000000000", "0100101110000000", "0100111011000000", "0101101011000000", "0101101010100000", "0101101010010000", "0101101010001000", "0101101101100000", "0101101100100000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101100111000", "0101101100110000", "0101101101100000", "0101101100101000", "0101101101001000", "0101000010000000", "0100110001000000", "0100111000000000", "0101000001000000", "0100101100000000", "0100110011000000", "0100110011000000", "0100110100000000", "0100110101000000", "0100110100000000", "0100110101000000", "0100110011000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100111000000000", "0100111110000000", "0101000000100000", "0100110100000000", "0100111000000000", "0100110111000000", "0100110011000000", "0100110001000000", "0100110001000000", "0100101110000000", "0100111110000000", "0101000100000000", "0101101111100000", "0101101111101000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101101101000", "0101101111101000", "0101101111101000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101110111000", "0101000100100000", "0101000111000000", "0101001000000000", "0101001000000000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000110000000", "0101000111000000", "0101000010100000", "0101000111000000", "0101000111100000", "0101001001000000", "0101001000100000", "0101000110100000", "0101000110100000", "0101000111100000", "0101000110000000", "0101000100100000", "0101000101000000", "0101000100100000", "0101000110100000", "0101000101000000", "0101000011000000", "0101000010000000", "0101000010100000", "0100111110000000", "0101000001100000", "0100111110000000", "0101000000000000", "0100110110000000", "0100110010000000", "0100110011000000", "0100111000000000", "0101101011101000", "0101101010100000", "0101101010010000", "0101101010001000", "0101101101100000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101101011000", "0101101100101000", "0101101100111000", "0101101101000000", "0101100010001000", "0100110011000000", "0100110010000000", "0100111101000000", "0100101000000000", "0100110010000000", "0100110011000000", "0100110101000000", "0100110110000000", "0100110100000000", "0100110101000000", "0100110100000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100111000000000", "0100111110000000", "0100111111000000", "0100110101000000", "0100110101000000", "0100110110000000", "0100110010000000", "0100110001000000", "0100110000000000", "0100101110000000", "0100111111000000", "0101000010000000", "0101101111101000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101110110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111101000", "0101101111011000", "0101101111111000", "0101101110011000", "0101000100000000", "0101000111000000", "0101000110000000", "0101000110100000", "0101000110100000", "0101000111000000", "0101000101100000", "0101000101100000", "0101000110100000", "0101000010000000", "0101000111000000", "0101000110100000", "0101001000000000", "0101000111100000", "0101000110000000", "0101000110100000", "0101000111100000", "0101000110000000", "0101000100100000", "0101000100100000", "0101000010100000", "0101000100100000", "0101000100000000", "0101000011100000", "0101000010000000", "0101000000100000", "0100110110000000", "0101000100100000", "0101000011100000", "0100110111000000", "0100110010000000", "0100110000000000", "0100110111000000", "0100110101000000", "0101101100001000", "0101101010100000", "0101101010010000", "0101101010000000", "0101101101100000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101101000000", "0101101101000000", "0101101100110000", "0101101101001000", "0101101100110000", "0101101101110000", "0100101100000000", "0100110010000000", "0100111100000000", "0100100000000000", "0100101110000000", "0100110010000000", "0100110110000000", "0100110111000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110011000000", "0100110100000000", "0100110111000000", "0100111010000000", "0100111111000000", "0100111110000000", "0100110101000000", "0100110100000000", "0100111000000000", "0100110100000000", "0100110001000000", "0100110000000000", "0100101110000000", "0100111101000000", "0100111110000000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111100000", "0101101111101000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101110001000", "0101000100000000", "0101001000100000", "0101000110100000", "0101000110100000", "0101000111000000", "0101000111100000", "0101000110100000", "0101000110000000", "0101000111000000", "0101000011100000", "0101000101100000", "0101000110100000", "0101000111100000", "0101000111100000", "0101000110100000", "0101000111100000", "0101000111100000", "0101000110000000", "0101000100100000", "0101000100000000", "0101000010000000", "0101000011100000", "0101000100000000", "0101000101000000", "0101000011000000", "0100111110000000", "0100110000000000", "0101000011000000", "0101000000000000", "0100110010000000", "0100101000000000", "0100110111000000", "0100110111000000", "0100110010000000", "0101101000010000", "0101101010100000", "0101101010010000", "0101101010000000", "0101101101100000", "0101101100101000", "0101101100110000", "0101101100110000", "0101101100111000", "0101101100110000", "0101101100111000", "0101101101000000", "0101101101001000", "0101101101011000", "0101101101001000", "0101101100110000", "0101101100110000", "0101101010010000", "0100110000000000", "0100101110000000", "0100111011000000", "0100100100000000", "0100101110000000", "0100110001000000", "0100110101000000", "0100110111000000", "0100110100000000", "0100110100000000", "0100110011000000", "0100110100000000", "0100110101000000", "0100110111000000", "0100111001000000", "0100111101000000", "0100111011000000", "0100110110000000", "0100110101000000", "0100111000000000", "0100110101000000", "0100110010000000", "0100110001000000", "0100110001000000", "0100111100000000", "0100110111000000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111101000", "0101101111010000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111100000", "0101101111100000", "0101101101011000", "0101000110000000", "0101001001100000", "0101000111000000", "0101000111100000", "0101001000000000", "0101000111000000", "0101000111000000", "0101000110100000", "0101000111100000", "0101000101100000", "0101000100000000", "0101000111100000", "0101000111100000", "0101000111000000", "0101000110100000", "0101000111100000", "0101000111000000", "0101000101000000", "0101000100100000", "0101000011100000", "0101000011100000", "0101000101000000", "0101000100000000", "0101000100100000", "0101000010000000", "0100111110000000", "0100110101000000", "0101000010000000", "0101000010000000", "0100110011000000", "0100110101000000", "0100110101000000", "0100110011000000", "0100110100000000", "0000000000000000", "0101101010100000", "0101101010010000", "0101101010001000", "0101101101100000", "0101101100101000", "0101101100110000", "0101101100111000", "0101101100111000", "0101101100110000", "0101101100111000", "0101101101000000", "0101101101001000", "0101101100101000", "0101101101000000", "0101101100100000", "0101101100110000", "0100110011000000", "0100101110000000", "0100110001000000", "0100110100000000", "0100101110000000", "0100110010000000", "0100110010000000", "0100110100000000", "0100110110000000", "0100110011000000", "0100110011000000", "0100110011000000", "0100110101000000", "0100110101000000", "0100110111000000", "0100110111000000", "0100111010000000", "0100111001000000", "0100110110000000", "0100110110000000", "0100110011000000", "0100110011000000", "0100110010000000", "0100110010000000", "0100110100000000", "0100111100000000", "0100110011000000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111010000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111110000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101101011000", "0101000101000000", "0101001000100000", "0101000111100000", "0101001000000000", "0101001000000000", "0101000101100000", "0101000110000000", "0101000101100000", "0101000111100000", "0101000110100000", "0101000011100000", "0101001000000000", "0101000111000000", "0101000110000000", "0101000110000000", "0101000111000000", "0101000101100000", "0101000100000000", "0101000011100000", "0101000011000000", "0101000101100000", "0101000111000000", "0101000011100000", "0101000010000000", "0100111110000000", "0100111101000000", "0100111101000000", "0101000010000000", "0100111010000000", "0100110011000000", "0100110000000000", "0100110011000000", "0100110100000000", "0100101000000000", "0100101100000000", "0101101010100000", "0101101010010000", "0101101010001000", "0101101101100000", "0101101100110000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101101000000", "0101101101000000", "0101101101000000", "0101101101001000", "0101101100100000", "0101101101000000", "0101101100111000", "0100110000000000", "0100110001000000", "0100101100000000", "0100110101000000", "0100111001000000", "0100101100000000", "0100110001000000", "0100110110000000", "0100110100000000", "0100110100000000", "0100110011000000", "0100110011000000", "0100110110000000", "0100110111000000", "0100110110000000", "0100111010000000", "0100111110000000", "0100110001000000", "0100111000000000", "0100110100000000", "0100110101000000", "0100110011000000", "0100110011000000", "0100101110000000", "0100110011000000", "0100111111000000", "0100111001000000", "0101101111111000", "0101101111101000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111100000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111100000", "0101101111111000", "0101101111011000", "0101101100001000", "0101000101100000", "0101001000100000", "0101001000100000", "0101001000100000", "0101000111100000", "0101000111100000", "0101000111000000", "0101000101000000", "0101001000000000", "0101000110000000", "0101000100000000", "0101000111100000", "0101001000000000", "0101001000000000", "0101001000000000", "0101000111100000", "0101000101100000", "0101000100100000", "0101000101000000", "0101000011000000", "0101000100100000", "0101000100100000", "0101000011100000", "0100111110000000", "0101000000100000", "0100111010000000", "0101000011000000", "0101000010000000", "0100110110000000", "0100101100000000", "0100110011000000", "0100110011000000", "0100100100000000", "0100011100000000", "0100100100000000", "0101101011001000", "0101101010100000", "0101101010010000", "0101101101101000", "0101101100110000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101101000000", "0101101101000000", "0101101101000000", "0101101100110000", "0101101101011000", "0101101100110000", "0101101010011000", "0100101110000000", "0100101010000000", "0100110100000000", "0100110001000000", "0100111010000000", "0100101110000000", "0100110010000000", "0100110111000000", "0100110101000000", "0100110101000000", "0100110100000000", "0100110100000000", "0100110100000000", "0100110110000000", "0100110100000000", "0100111001000000", "0100111100000000", "0100101110000000", "0100110111000000", "0100110011000000", "0100110100000000", "0100110011000000", "0100110010000000", "0100110000000000", "0100110100000000", "0101000000000000", "0100111110000000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101110111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111101000", "0101101111111000", "0101101111011000", "0101101111011000", "0101101001000000", "0101000100100000", "0101001001100000", "0101000111000000", "0101000111100000", "0101000111000000", "0101001000000000", "0101001000000000", "0101000110000000", "0101001000000000", "0101000101100000", "0101000011100000", "0101000111000000", "0101000111000000", "0101000110100000", "0101000110100000", "0101000111000000", "0101000101100000", "0101000100000000", "0101000100100000", "0101000011000000", "0101000001000000", "0101000101000000", "0101000100000000", "0100111101000000", "0100111100000000", "0100110000000000", "0101000010100000", "0100111111000000", "0100110100000000", "0100110100000000", "0100111010000000", "0100110100000000", "0100101010000000", "0100100110000000", "0100100010000000", "0101101010111000", "0101101010010000", "0101101010001000", "0101101101101000", "0101101100111000", "0101101101000000", "0101101101000000", "0101101100111000", "0101101100111000", "0101101100111000", "0101101101000000", "0101101101001000", "0101101101010000", "0101101100100000", "0101101100111000", "0101000001000000", "0100101110000000", "0100110001000000", "0100101100000000", "0100110010000000", "0100111001000000", "0100101110000000", "0100110010000000", "0100110111000000", "0100110101000000", "0100110100000000", "0100110100000000", "0100110100000000", "0100110100000000", "0100110110000000", "0100110100000000", "0100111000000000", "0100111011000000", "0100101100000000", "0100110111000000", "0100110100000000", "0100110100000000", "0100110011000000", "0100110001000000", "0100110001000000", "0100110100000000", "0101000000000000", "0101000010100000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101110001000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111101000", "0101101110110000", "0101011010010000", "0101000111000000", "0101001001100000", "0101001000000000", "0101000111000000", "0101000111000000", "0101001000000000", "0101001000100000", "0101000110000000", "0101001000000000", "0101000110000000", "0101000100000000", "0101000110100000", "0101000110100000", "0101000110000000", "0101000110000000", "0101000110000000", "0101000101000000", "0101000100000000", "0101000100000000", "0101000010100000", "0101000001000000", "0101000101000000", "0101000100000000", "0100111011000000", "0100111000000000", "0100110000000000", "0101000010100000", "0100111100000000", "0100110100000000", "0100111000000000", "0100111010000000", "0100110001000000", "0100101110000000", "0100110011000000", "0100110001000000", "0101101010110000", "0101101010001000", "0101101010000000", "0101101101100000", "0101101101000000", "0101101101000000", "0101101101000000", "0101101100111000", "0101101100111000", "0101101101000000", "0101101101000000", "0101101101000000", "0101101101001000", "0101101101000000", "0101101100100000", "0100100010000000", "0100110000000000", "0100101000000000", "0100101110000000", "0100110100000000", "0100111000000000", "0100101100000000", "0100110000000000", "0100110101000000", "0100110100000000", "0100110011000000", "0100110011000000", "0100110011000000", "0100110101000000", "0100110111000000", "0100110101000000", "0100111001000000", "0100111011000000", "0100101100000000", "0100111000000000", "0100110101000000", "0100110101000000", "0100110101000000", "0100110010000000", "0100110001000000", "0100110100000000", "0101000000000000", "0101000100100000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101101100000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111110000", "0101101111111000", "0101101111111000", "0101101111110000", "0101101111111000", "0101101111011000", "0101101111111000", "0101101110100000", "0100110111000000", "0101001001000000", "0101001010000000", "0101001000100000", "0101000111100000", "0101000111000000", "0101001000000000", "0101001000000000", "0101000101100000", "0101000111100000", "0101000110100000", "0101000110000000", "0101000111000000", "0101000111000000", "0101000110000000", "0101000110000000", "0101000110100000", "0101000101000000", "0101000011100000", "0101000011000000", "0101000001000000", "0101000100000000", "0101000100000000", "0101000011000000", "0100111001000000", "0100110110000000", "0100111010000000", "0101000010100000", "0100111000000000", "0100110110000000", "0100111010000000", "0100110110000000", "0100101110000000", "0100110010000000", "0100111000000000", "0100111001000000", "0101101010111000", "0101101010010000", "0101101010000000", "0101101101100000"
	);
	
	--signal tmp : std_logic := '0';
	--signal i,j : integer := 0;
begin
	conv_dut  : conv2d generic map (100, 100, 7, 7) port map (clk, img_rom, log_rom, filtered_img);
	
--	process (clk)
--	begin
--		if (rising_edge(clk)) then
--			for i in 0 to 4 loop
--				for j in 0 to 4 loop
--						--tmp <= not tmp;
--						report ("i and j are " & integer'image(i) & " " & integer'image(j));
--				end loop;
--			end loop;
--		end if;
--	end process;
	
--	process (clk)
--	begin
--		if (rising_edge(clk)) then
--			if (i < 3) then
--				if (j < 3) then
--					report ("i and j are " & integer'image(i) & " " & integer'image(j));
--					j <= j+1;
--				end if;
--				if (j = 3-1) then
--					j <= 0;
--					i <= i + 1;
--				end if;
--			end if;
--		end if;
--	end process;
	
end architecture;